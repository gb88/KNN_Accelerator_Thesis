// nios_sys.v

// Generated using ACDS version 12.1 177 at 2014.07.10.19:46:42

`timescale 1 ps / 1 ps
module nios_sys (
		output wire        altpll_0_c1_clk,                         //                 altpll_0_c1.clk
		output wire        FIFO_wr_n_from_the_usbFIFOCtrl_0,        //   usbFIFOCtrl_0_conduit_end.export
		input  wire        reset_n,                                 //          clk_0_clk_in_reset.reset_n
		output wire [11:0] zs_addr_from_the_sdram_0,                //                sdram_0_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram_0,                  //                            .ba
		output wire        zs_cas_n_from_the_sdram_0,               //                            .cas_n
		output wire        zs_cke_from_the_sdram_0,                 //                            .cke
		output wire        zs_cs_n_from_the_sdram_0,                //                            .cs_n
		inout  wire [31:0] zs_dq_to_and_from_the_sdram_0,           //                            .dq
		output wire [3:0]  zs_dqm_from_the_sdram_0,                 //                            .dqm
		output wire        zs_ras_n_from_the_sdram_0,               //                            .ras_n
		output wire        zs_we_n_from_the_sdram_0,                //                            .we_n
		output wire [7:0]  out_port_from_the_pio_0,                 //   pio_0_external_connection.export
		output wire [2:0]  led_from_the_usbFIFOCtrl_0,              // usbFIFOCtrl_0_conduit_end_8.export
		input  wire        FLAGC_n_to_the_usbFIFOCtrl_0,            // usbFIFOCtrl_0_conduit_end_7.export
		input  wire        FLAGB_n_to_the_usbFIFOCtrl_0,            // usbFIFOCtrl_0_conduit_end_6.export
		inout  wire [15:0] FIFO_data_to_and_from_the_usbFIFOCtrl_0, // usbFIFOCtrl_0_conduit_end_5.export
		output wire [1:0]  FIFO_add_from_the_usbFIFOCtrl_0,         // usbFIFOCtrl_0_conduit_end_4.export
		input  wire        clk_1_clk_in_clk,                        //                clk_1_clk_in.clk
		output wire        FIFO_pktend_from_the_usbFIFOCtrl_0,      // usbFIFOCtrl_0_conduit_end_3.export
		output wire        FIFO_oe_n_from_the_usbFIFOCtrl_0,        // usbFIFOCtrl_0_conduit_end_2.export
		output wire        FIFO_rd_n_from_the_usbFIFOCtrl_0,        // usbFIFOCtrl_0_conduit_end_1.export
		input  wire        clk_0,                                   //                clk_0_clk_in.clk
		input  wire        clk_1_clk_in_reset_reset_n               //          clk_1_clk_in_reset.reset_n
	);

	wire   [15:0] distancecore_0_dist_export;                                                                               // distancecore_0:Dist -> knnclasscore:Dist0
	wire   [15:0] distancecore_1_dist_export;                                                                               // distancecore_1:Dist -> knnclasscore:Dist1
	wire          distancecore_0_endcomp_export;                                                                            // distancecore_0:EndComp -> knnclasscore:EndComp0
	wire          distancecore_1_endcomp_export;                                                                            // distancecore_1:EndComp -> knnclasscore:EndComp1
	wire          knnclasscore_go0_export;                                                                                  // knnclasscore:Go0 -> distancecore_0:Go
	wire          knnclasscore_go1_export;                                                                                  // knnclasscore:Go1 -> distancecore_1:Go
	wire    [3:0] distancecore_0_cl_export;                                                                                 // distancecore_0:Cl -> knnclasscore:Cl0
	wire    [3:0] distancecore_1_cl_export;                                                                                 // distancecore_1:Cl -> knnclasscore:Cl1
	wire    [7:0] ndimreg_ndim0_export;                                                                                     // NDimReg:NDim0 -> distancecore_0:NDim
	wire    [7:0] ndimreg_ndim1_export;                                                                                     // NDimReg:NDim1 -> distancecore_1:NDim
	wire    [7:0] ntrreg_0_ntr_export;                                                                                      // NTrReg_0:NTr -> distancecore_0:NTr
	wire    [7:0] ntrreg_1_ntr_export;                                                                                      // NTrReg_1:NTr -> distancecore_1:NTr
	wire          fullreg_1_full_export;                                                                                    // FullReg_1:Full -> distancecore_1:Full
	wire          fullreg_0_full_export;                                                                                    // FullReg_0:Full -> distancecore_0:Full
	wire          distancecore_0_empty_export;                                                                              // distancecore_0:Empty -> emptyreg_0:Empty
	wire          distancecore_1_empty_export;                                                                              // distancecore_1:Empty -> emptyreg_1:Empty
	wire          distancecore_0_endtsetout_export;                                                                         // distancecore_0:EndTSetOut -> knnclasscore:EndTSet0
	wire          distancecore_1_endtsetout_export;                                                                         // distancecore_1:EndTSetOut -> knnclasscore:EndTSet1
	wire          endtsetreg_0_endtset_export;                                                                              // EndTSetReg_0:EndTSet -> distancecore_0:EndTSetIn
	wire          endtsetreg_1_endtset_export;                                                                              // EndTSetReg_1:EndTSet -> distancecore_1:EndTSetIn
	wire          knnclasscore_distreset0_export;                                                                           // knnclasscore:DistReset0 -> distancecore_0:reset
	wire          knnclasscore_distreset1_export;                                                                           // knnclasscore:DistReset1 -> distancecore_1:reset
	wire          knnclasscore_drop1_export;                                                                                // knnclasscore:Drop1 -> distancecore_1:Drop
	wire          knnclasscore_drop0_export;                                                                                // knnclasscore:Drop0 -> distancecore_0:Drop
	wire   [15:0] baseqaddr_0_qaddress0_export;                                                                             // baseqaddr_0:QAddress0 -> distancecore_0:QAddress
	wire   [15:0] baseqaddr_0_qaddress1_export;                                                                             // baseqaddr_0:QAddress1 -> distancecore_1:QAddress
	wire          altpll_0_c2_clk;                                                                                          // altpll_0:c2 -> [addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, cache_0:clk, cache_0:clk2, cache_0_s1_translator:clk, cache_0_s1_translator_avalon_universal_slave_0_agent:clk, cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cache_0_s2_translator:clk, cache_0_s2_translator_avalon_universal_slave_0_agent:clk, cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cache_1:clk, cache_1:clk2, cache_1_s1_translator:clk, cache_1_s1_translator_avalon_universal_slave_0_agent:clk, cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cache_1_s2_translator:clk, cache_1_s2_translator_avalon_universal_slave_0_agent:clk, cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cache_2:clk, cache_2:clk2, cache_2_s1_translator:clk, cache_2_s1_translator_avalon_universal_slave_0_agent:clk, cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cache_2_s2_translator:clk, cache_2_s2_translator_avalon_universal_slave_0_agent:clk, cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_005:clk, cmd_xbar_mux_023:clk, cmd_xbar_mux_024:clk, cmd_xbar_mux_025:clk, cpu_0:clk, cpu_0_data_master_translator:clk, cpu_0_data_master_translator_avalon_universal_master_0_agent:clk, cpu_0_instruction_master_translator:clk, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:clk, crosser:in_clk, crosser_001:in_clk, crosser_002:in_clk, crosser_003:in_clk, crosser_004:in_clk, crosser_005:in_clk, crosser_006:in_clk, crosser_007:in_clk, crosser_008:in_clk, crosser_009:in_clk, crosser_010:in_clk, crosser_011:in_clk, crosser_012:in_clk, crosser_013:in_clk, crosser_014:in_clk, crosser_015:in_clk, crosser_016:in_clk, crosser_017:out_clk, crosser_018:out_clk, crosser_019:out_clk, crosser_020:out_clk, crosser_021:out_clk, crosser_022:out_clk, crosser_023:out_clk, crosser_024:out_clk, crosser_025:out_clk, crosser_026:out_clk, crosser_027:out_clk, crosser_028:out_clk, crosser_029:out_clk, crosser_030:out_clk, crosser_031:out_clk, crosser_032:out_clk, crosser_033:out_clk, crosser_034:out_clk, crosser_035:out_clk, crosser_036:out_clk, crosser_037:in_clk, crosser_038:in_clk, crosser_039:in_clk, crosser_040:out_clk, crosser_041:in_clk, crosser_042:out_clk, crosser_043:in_clk, crosser_044:out_clk, crosser_045:in_clk, dma:clk, dma_control_port_slave_translator:clk, dma_control_port_slave_translator_avalon_universal_slave_0_agent:clk, dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dma_read_master_translator:clk, dma_read_master_translator_avalon_universal_master_0_agent:clk, dma_write_master_translator:clk, dma_write_master_translator_avalon_universal_master_0_agent:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_005:clk, id_router_006:clk, id_router_023:clk, id_router_024:clk, id_router_025:clk, id_router_026:clk, id_router_027:clk, id_router_028:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, performance_counter_0:clk, performance_counter_0_control_slave_translator:clk, performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:clk, performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_0:clk, pio_0_s1_translator:clk, pio_0_s1_translator_avalon_universal_slave_0_agent:clk, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_023:clk, rsp_xbar_demux_024:clk, rsp_xbar_demux_025:clk, rsp_xbar_demux_026:clk, rsp_xbar_demux_027:clk, rsp_xbar_demux_028:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rsp_xbar_mux_003:clk, rst_controller:clk, sdram_controller:clk, sdram_controller_s1_translator:clk, sdram_controller_s1_translator_avalon_universal_slave_0_agent:clk, sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire   [15:0] skipaddrreg_0_skipaddr0_export;                                                                           // skipaddrreg_0:SkipAddr0 -> distancecore_0:SkipAddr
	wire   [15:0] skipaddrreg_0_skipaddr1_export;                                                                           // skipaddrreg_0:SkipAddr1 -> distancecore_1:SkipAddr
	wire          altpll_0_c0_clk;                                                                                          // altpll_0:c0 -> [burst_adapter:clk, crosser:out_clk, crosser_017:in_clk, id_router_004:clk, rsp_xbar_demux_004:clk, rst_controller_001:clk, usbFIFOCtrl_0:clk, usbFIFOCtrl_0_avalon_slave_0_translator:clk, usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk]
	wire          altpll_1_c0_clk;                                                                                          // altpll_1:c0 -> [EndTSetReg_0:clk, EndTSetReg_0_avalon_slave_0_translator:clk, EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, EndTSetReg_1:clk, EndTSetReg_1_avalon_slave_0_translator:clk, EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, EndTSetReg_2:clk, EndTSetReg_2_avalon_slave_0_translator:clk, EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FullReg_0:clk, FullReg_0_avalon_slave_0_translator:clk, FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FullReg_1:clk, FullReg_1_avalon_slave_0_translator:clk, FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, FullReg_2:clk, FullReg_2_avalon_slave_0_translator:clk, FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, NDimReg:clk, NDimReg_avalon_slave_0_translator:clk, NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, NTrReg_0:clk, NTrReg_0_avalon_slave_0_translator:clk, NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, NTrReg_1:clk, NTrReg_1_avalon_slave_0_translator:clk, NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, NTrReg_2:clk, NTrReg_2_avalon_slave_0_translator:clk, NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router_004:clk, addr_router_005:clk, addr_router_006:clk, addr_router_007:clk, addr_router_008:clk, addr_router_009:clk, baseqaddr_0:clk, baseqaddr_0_avalon_slave_0_translator:clk, baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux_004:clk, cmd_xbar_demux_005:clk, cmd_xbar_demux_006:clk, cmd_xbar_demux_007:clk, cmd_xbar_demux_008:clk, cmd_xbar_demux_009:clk, crosser_001:out_clk, crosser_002:out_clk, crosser_003:out_clk, crosser_004:out_clk, crosser_005:out_clk, crosser_006:out_clk, crosser_007:out_clk, crosser_008:out_clk, crosser_009:out_clk, crosser_010:out_clk, crosser_011:out_clk, crosser_012:out_clk, crosser_013:out_clk, crosser_014:out_clk, crosser_015:out_clk, crosser_016:out_clk, crosser_018:in_clk, crosser_019:in_clk, crosser_020:in_clk, crosser_021:in_clk, crosser_022:in_clk, crosser_023:in_clk, crosser_024:in_clk, crosser_025:in_clk, crosser_026:in_clk, crosser_027:in_clk, crosser_028:in_clk, crosser_029:in_clk, crosser_030:in_clk, crosser_031:in_clk, crosser_032:in_clk, crosser_033:in_clk, crosser_034:in_clk, crosser_035:in_clk, crosser_036:in_clk, crosser_037:out_clk, crosser_038:out_clk, crosser_039:out_clk, crosser_040:in_clk, crosser_041:out_clk, crosser_042:in_clk, crosser_043:out_clk, crosser_044:in_clk, crosser_045:out_clk, distancecore_0:Clk, distancecore_0_avalon_master_1_translator:clk, distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:clk, distancecore_0_avalon_master_translator:clk, distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:clk, distancecore_1:Clk, distancecore_1_avalon_master_1_translator:clk, distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:clk, distancecore_1_avalon_master_translator:clk, distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:clk, distancecore_2:Clk, distancecore_2_avalon_master_1_translator:clk, distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:clk, distancecore_2_avalon_master_translator:clk, distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:clk, emptyreg_0:clk, emptyreg_0_avalon_slave_0_translator:clk, emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, emptyreg_1:clk, emptyreg_1_avalon_slave_0_translator:clk, emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, emptyreg_2:clk, emptyreg_2_avalon_slave_0_translator:clk, emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, id_router_019:clk, id_router_020:clk, id_router_021:clk, id_router_022:clk, knnclasscore:Clk, knnclasscore_avalon_slave_0_translator:clk, knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_demux_019:clk, rsp_xbar_demux_020:clk, rsp_xbar_demux_021:clk, rsp_xbar_demux_022:clk, rst_controller_003:clk, skipaddrreg_0:clk, skipaddrreg_0_avalon_slave_0_translator:clk, skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire          distancecore_0_overflow_export;                                                                           // distancecore_0:Overflow -> knnclasscore:Overflow0
	wire          distancecore_1_overflow_export;                                                                           // distancecore_1:Overflow -> knnclasscore:Overflow1
	wire   [15:0] baseqaddr_0_qaddress2_export;                                                                             // baseqaddr_0:QAddress2 -> distancecore_2:QAddress
	wire          distancecore_2_empty_export;                                                                              // distancecore_2:Empty -> emptyreg_2:Empty
	wire          endtsetreg_2_endtset_export;                                                                              // EndTSetReg_2:EndTSet -> distancecore_2:EndTSetIn
	wire          fullreg_2_full_export;                                                                                    // FullReg_2:Full -> distancecore_2:Full
	wire    [7:0] ndimreg_ndim2_export;                                                                                     // NDimReg:NDim2 -> distancecore_2:NDim
	wire    [7:0] ntrreg_2_ntr_export;                                                                                      // NTrReg_2:NTr -> distancecore_2:NTr
	wire   [15:0] skipaddrreg_0_skipaddr2_export;                                                                           // skipaddrreg_0:SkipAddr2 -> distancecore_2:SkipAddr
	wire          knnclasscore_drop2_export;                                                                                // knnclasscore:Drop2 -> distancecore_2:Drop
	wire          knnclasscore_distreset2_export;                                                                           // knnclasscore:DistReset2 -> distancecore_2:reset
	wire   [15:0] distancecore_2_dist_export;                                                                               // distancecore_2:Dist -> knnclasscore:Dist2
	wire          distancecore_2_endtsetout_export;                                                                         // distancecore_2:EndTSetOut -> knnclasscore:EndTSet2
	wire    [3:0] distancecore_2_cl_export;                                                                                 // distancecore_2:Cl -> knnclasscore:Cl2
	wire          distancecore_2_endcomp_export;                                                                            // distancecore_2:EndComp -> knnclasscore:EndComp2
	wire          knnclasscore_go2_export;                                                                                  // knnclasscore:Go2 -> distancecore_2:Go
	wire          distancecore_2_overflow_export;                                                                           // distancecore_2:Overflow -> knnclasscore:Overflow2
	wire          cpu_0_instruction_master_waitrequest;                                                                     // cpu_0_instruction_master_translator:av_waitrequest -> cpu_0:i_waitrequest
	wire   [25:0] cpu_0_instruction_master_address;                                                                         // cpu_0:i_address -> cpu_0_instruction_master_translator:av_address
	wire          cpu_0_instruction_master_read;                                                                            // cpu_0:i_read -> cpu_0_instruction_master_translator:av_read
	wire   [31:0] cpu_0_instruction_master_readdata;                                                                        // cpu_0_instruction_master_translator:av_readdata -> cpu_0:i_readdata
	wire          cpu_0_data_master_waitrequest;                                                                            // cpu_0_data_master_translator:av_waitrequest -> cpu_0:d_waitrequest
	wire   [31:0] cpu_0_data_master_writedata;                                                                              // cpu_0:d_writedata -> cpu_0_data_master_translator:av_writedata
	wire   [25:0] cpu_0_data_master_address;                                                                                // cpu_0:d_address -> cpu_0_data_master_translator:av_address
	wire          cpu_0_data_master_write;                                                                                  // cpu_0:d_write -> cpu_0_data_master_translator:av_write
	wire          cpu_0_data_master_read;                                                                                   // cpu_0:d_read -> cpu_0_data_master_translator:av_read
	wire   [31:0] cpu_0_data_master_readdata;                                                                               // cpu_0_data_master_translator:av_readdata -> cpu_0:d_readdata
	wire    [3:0] cpu_0_data_master_byteenable;                                                                             // cpu_0:d_byteenable -> cpu_0_data_master_translator:av_byteenable
	wire          dma_read_master_waitrequest;                                                                              // dma_read_master_translator:av_waitrequest -> dma:read_waitrequest
	wire   [24:0] dma_read_master_address;                                                                                  // dma:read_address -> dma_read_master_translator:av_address
	wire          dma_read_master_chipselect;                                                                               // dma:read_chipselect -> dma_read_master_translator:av_chipselect
	wire          dma_read_master_read;                                                                                     // dma:read_read_n -> dma_read_master_translator:av_read
	wire   [31:0] dma_read_master_readdata;                                                                                 // dma_read_master_translator:av_readdata -> dma:read_readdata
	wire          dma_read_master_readdatavalid;                                                                            // dma_read_master_translator:av_readdatavalid -> dma:read_readdatavalid
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                             // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire   [11:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                               // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                            // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                 // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                 // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                              // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                            // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire   [31:0] dma_control_port_slave_translator_avalon_anti_slave_0_writedata;                                          // dma_control_port_slave_translator:av_writedata -> dma:dma_ctl_writedata
	wire    [2:0] dma_control_port_slave_translator_avalon_anti_slave_0_address;                                            // dma_control_port_slave_translator:av_address -> dma:dma_ctl_address
	wire          dma_control_port_slave_translator_avalon_anti_slave_0_chipselect;                                         // dma_control_port_slave_translator:av_chipselect -> dma:dma_ctl_chipselect
	wire          dma_control_port_slave_translator_avalon_anti_slave_0_write;                                              // dma_control_port_slave_translator:av_write -> dma:dma_ctl_write_n
	wire   [31:0] dma_control_port_slave_translator_avalon_anti_slave_0_readdata;                                           // dma:dma_ctl_readdata -> dma_control_port_slave_translator:av_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                 // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                     // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                       // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                        // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                    // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] pio_0_s1_translator_avalon_anti_slave_0_writedata;                                                        // pio_0_s1_translator:av_writedata -> pio_0:writedata
	wire    [1:0] pio_0_s1_translator_avalon_anti_slave_0_address;                                                          // pio_0_s1_translator:av_address -> pio_0:address
	wire          pio_0_s1_translator_avalon_anti_slave_0_chipselect;                                                       // pio_0_s1_translator:av_chipselect -> pio_0:chipselect
	wire          pio_0_s1_translator_avalon_anti_slave_0_write;                                                            // pio_0_s1_translator:av_write -> pio_0:write_n
	wire   [31:0] pio_0_s1_translator_avalon_anti_slave_0_readdata;                                                         // pio_0:readdata -> pio_0_s1_translator:av_readdata
	wire   [15:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                    // usbFIFOCtrl_0_avalon_slave_0_translator:av_writedata -> usbFIFOCtrl_0:writedata
	wire    [1:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                      // usbFIFOCtrl_0_avalon_slave_0_translator:av_address -> usbFIFOCtrl_0:address
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                   // usbFIFOCtrl_0_avalon_slave_0_translator:av_chipselect -> usbFIFOCtrl_0:chipselect
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                        // usbFIFOCtrl_0_avalon_slave_0_translator:av_write -> usbFIFOCtrl_0:write
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                         // usbFIFOCtrl_0_avalon_slave_0_translator:av_read -> usbFIFOCtrl_0:read
	wire   [15:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                     // usbFIFOCtrl_0:readdata -> usbFIFOCtrl_0_avalon_slave_0_translator:av_readdata
	wire    [1:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                                   // usbFIFOCtrl_0_avalon_slave_0_translator:av_byteenable -> usbFIFOCtrl_0:byteenable
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest;                                           // sdram_controller:za_waitrequest -> sdram_controller_s1_translator:av_waitrequest
	wire   [31:0] sdram_controller_s1_translator_avalon_anti_slave_0_writedata;                                             // sdram_controller_s1_translator:av_writedata -> sdram_controller:az_data
	wire   [22:0] sdram_controller_s1_translator_avalon_anti_slave_0_address;                                               // sdram_controller_s1_translator:av_address -> sdram_controller:az_addr
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_chipselect;                                            // sdram_controller_s1_translator:av_chipselect -> sdram_controller:az_cs
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_write;                                                 // sdram_controller_s1_translator:av_write -> sdram_controller:az_wr_n
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_read;                                                  // sdram_controller_s1_translator:av_read -> sdram_controller:az_rd_n
	wire   [31:0] sdram_controller_s1_translator_avalon_anti_slave_0_readdata;                                              // sdram_controller:za_data -> sdram_controller_s1_translator:av_readdata
	wire          sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid;                                         // sdram_controller:za_valid -> sdram_controller_s1_translator:av_readdatavalid
	wire    [3:0] sdram_controller_s1_translator_avalon_anti_slave_0_byteenable;                                            // sdram_controller_s1_translator:av_byteenable -> sdram_controller:az_be_n
	wire   [31:0] performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata;                             // performance_counter_0_control_slave_translator:av_writedata -> performance_counter_0:writedata
	wire    [3:0] performance_counter_0_control_slave_translator_avalon_anti_slave_0_address;                               // performance_counter_0_control_slave_translator:av_address -> performance_counter_0:address
	wire          performance_counter_0_control_slave_translator_avalon_anti_slave_0_write;                                 // performance_counter_0_control_slave_translator:av_write -> performance_counter_0:write
	wire   [31:0] performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata;                              // performance_counter_0:readdata -> performance_counter_0_control_slave_translator:av_readdata
	wire          performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer;                         // performance_counter_0_control_slave_translator:av_begintransfer -> performance_counter_0:begintransfer
	wire   [31:0] ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                          // NDimReg_avalon_slave_0_translator:av_writedata -> NDimReg:writedata
	wire    [1:0] ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_address;                                            // NDimReg_avalon_slave_0_translator:av_address -> NDimReg:address
	wire          ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                         // NDimReg_avalon_slave_0_translator:av_chipselect -> NDimReg:chipselect
	wire          ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_write;                                              // NDimReg_avalon_slave_0_translator:av_write -> NDimReg:write
	wire          ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_read;                                               // NDimReg_avalon_slave_0_translator:av_read -> NDimReg:read
	wire   [31:0] ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                           // NDimReg:readdata -> NDimReg_avalon_slave_0_translator:av_readdata
	wire   [31:0] endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                     // EndTSetReg_0_avalon_slave_0_translator:av_writedata -> EndTSetReg_0:writedata
	wire    [1:0] endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                       // EndTSetReg_0_avalon_slave_0_translator:av_address -> EndTSetReg_0:address
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                    // EndTSetReg_0_avalon_slave_0_translator:av_chipselect -> EndTSetReg_0:chipselect
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                         // EndTSetReg_0_avalon_slave_0_translator:av_write -> EndTSetReg_0:write
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                          // EndTSetReg_0_avalon_slave_0_translator:av_read -> EndTSetReg_0:read
	wire   [31:0] endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                      // EndTSetReg_0:readdata -> EndTSetReg_0_avalon_slave_0_translator:av_readdata
	wire   [31:0] fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                        // FullReg_0_avalon_slave_0_translator:av_writedata -> FullReg_0:writedata
	wire    [1:0] fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                          // FullReg_0_avalon_slave_0_translator:av_address -> FullReg_0:address
	wire          fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                       // FullReg_0_avalon_slave_0_translator:av_chipselect -> FullReg_0:chipselect
	wire          fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                            // FullReg_0_avalon_slave_0_translator:av_write -> FullReg_0:write
	wire          fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                             // FullReg_0_avalon_slave_0_translator:av_read -> FullReg_0:read
	wire   [31:0] fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                         // FullReg_0:readdata -> FullReg_0_avalon_slave_0_translator:av_readdata
	wire   [31:0] fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                        // FullReg_1_avalon_slave_0_translator:av_writedata -> FullReg_1:writedata
	wire    [1:0] fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address;                                          // FullReg_1_avalon_slave_0_translator:av_address -> FullReg_1:address
	wire          fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                       // FullReg_1_avalon_slave_0_translator:av_chipselect -> FullReg_1:chipselect
	wire          fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write;                                            // FullReg_1_avalon_slave_0_translator:av_write -> FullReg_1:write
	wire          fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read;                                             // FullReg_1_avalon_slave_0_translator:av_read -> FullReg_1:read
	wire   [31:0] fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                         // FullReg_1:readdata -> FullReg_1_avalon_slave_0_translator:av_readdata
	wire   [31:0] ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                         // NTrReg_0_avalon_slave_0_translator:av_writedata -> NTrReg_0:writedata
	wire    [1:0] ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                           // NTrReg_0_avalon_slave_0_translator:av_address -> NTrReg_0:address
	wire          ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                        // NTrReg_0_avalon_slave_0_translator:av_chipselect -> NTrReg_0:chipselect
	wire          ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                             // NTrReg_0_avalon_slave_0_translator:av_write -> NTrReg_0:write
	wire          ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                              // NTrReg_0_avalon_slave_0_translator:av_read -> NTrReg_0:read
	wire   [31:0] ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                          // NTrReg_0:readdata -> NTrReg_0_avalon_slave_0_translator:av_readdata
	wire   [31:0] ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                         // NTrReg_1_avalon_slave_0_translator:av_writedata -> NTrReg_1:writedata
	wire    [1:0] ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address;                                           // NTrReg_1_avalon_slave_0_translator:av_address -> NTrReg_1:address
	wire          ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                        // NTrReg_1_avalon_slave_0_translator:av_chipselect -> NTrReg_1:chipselect
	wire          ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write;                                             // NTrReg_1_avalon_slave_0_translator:av_write -> NTrReg_1:write
	wire          ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read;                                              // NTrReg_1_avalon_slave_0_translator:av_read -> NTrReg_1:read
	wire   [31:0] ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                          // NTrReg_1:readdata -> NTrReg_1_avalon_slave_0_translator:av_readdata
	wire   [31:0] emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                       // emptyreg_0_avalon_slave_0_translator:av_writedata -> emptyreg_0:writedata
	wire    [1:0] emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                         // emptyreg_0_avalon_slave_0_translator:av_address -> emptyreg_0:address
	wire          emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                      // emptyreg_0_avalon_slave_0_translator:av_chipselect -> emptyreg_0:chipselect
	wire          emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                           // emptyreg_0_avalon_slave_0_translator:av_write -> emptyreg_0:write
	wire          emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                            // emptyreg_0_avalon_slave_0_translator:av_read -> emptyreg_0:read
	wire   [31:0] emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                        // emptyreg_0:readdata -> emptyreg_0_avalon_slave_0_translator:av_readdata
	wire   [31:0] emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                       // emptyreg_1_avalon_slave_0_translator:av_writedata -> emptyreg_1:writedata
	wire    [1:0] emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address;                                         // emptyreg_1_avalon_slave_0_translator:av_address -> emptyreg_1:address
	wire          emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                      // emptyreg_1_avalon_slave_0_translator:av_chipselect -> emptyreg_1:chipselect
	wire          emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write;                                           // emptyreg_1_avalon_slave_0_translator:av_write -> emptyreg_1:write
	wire          emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read;                                            // emptyreg_1_avalon_slave_0_translator:av_read -> emptyreg_1:read
	wire   [31:0] emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                        // emptyreg_1:readdata -> emptyreg_1_avalon_slave_0_translator:av_readdata
	wire   [31:0] endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                     // EndTSetReg_1_avalon_slave_0_translator:av_writedata -> EndTSetReg_1:writedata
	wire    [1:0] endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address;                                       // EndTSetReg_1_avalon_slave_0_translator:av_address -> EndTSetReg_1:address
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                    // EndTSetReg_1_avalon_slave_0_translator:av_chipselect -> EndTSetReg_1:chipselect
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write;                                         // EndTSetReg_1_avalon_slave_0_translator:av_write -> EndTSetReg_1:write
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read;                                          // EndTSetReg_1_avalon_slave_0_translator:av_read -> EndTSetReg_1:read
	wire   [31:0] endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                      // EndTSetReg_1:readdata -> EndTSetReg_1_avalon_slave_0_translator:av_readdata
	wire   [31:0] baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                      // baseqaddr_0_avalon_slave_0_translator:av_writedata -> baseqaddr_0:writedata
	wire    [1:0] baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                        // baseqaddr_0_avalon_slave_0_translator:av_address -> baseqaddr_0:address
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                     // baseqaddr_0_avalon_slave_0_translator:av_chipselect -> baseqaddr_0:chipselect
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                          // baseqaddr_0_avalon_slave_0_translator:av_write -> baseqaddr_0:write
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                           // baseqaddr_0_avalon_slave_0_translator:av_read -> baseqaddr_0:read
	wire   [31:0] baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                       // baseqaddr_0:readdata -> baseqaddr_0_avalon_slave_0_translator:av_readdata
	wire   [31:0] skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                    // skipaddrreg_0_avalon_slave_0_translator:av_writedata -> skipaddrreg_0:writedata
	wire    [1:0] skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                      // skipaddrreg_0_avalon_slave_0_translator:av_address -> skipaddrreg_0:address
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                   // skipaddrreg_0_avalon_slave_0_translator:av_chipselect -> skipaddrreg_0:chipselect
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                        // skipaddrreg_0_avalon_slave_0_translator:av_write -> skipaddrreg_0:write
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                         // skipaddrreg_0_avalon_slave_0_translator:av_read -> skipaddrreg_0:read
	wire   [31:0] skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                     // skipaddrreg_0:readdata -> skipaddrreg_0_avalon_slave_0_translator:av_readdata
	wire   [31:0] knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                     // knnclasscore_avalon_slave_0_translator:av_writedata -> knnclasscore:writedata
	wire    [4:0] knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_address;                                       // knnclasscore_avalon_slave_0_translator:av_address -> knnclasscore:address
	wire          knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                    // knnclasscore_avalon_slave_0_translator:av_chipselect -> knnclasscore:chipselect
	wire          knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_write;                                         // knnclasscore_avalon_slave_0_translator:av_write -> knnclasscore:write
	wire          knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_read;                                          // knnclasscore_avalon_slave_0_translator:av_read -> knnclasscore:read
	wire   [31:0] knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                      // knnclasscore:readdata -> knnclasscore_avalon_slave_0_translator:av_readdata
	wire   [31:0] emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                       // emptyreg_2_avalon_slave_0_translator:av_writedata -> emptyreg_2:writedata
	wire    [1:0] emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address;                                         // emptyreg_2_avalon_slave_0_translator:av_address -> emptyreg_2:address
	wire          emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                      // emptyreg_2_avalon_slave_0_translator:av_chipselect -> emptyreg_2:chipselect
	wire          emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write;                                           // emptyreg_2_avalon_slave_0_translator:av_write -> emptyreg_2:write
	wire          emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read;                                            // emptyreg_2_avalon_slave_0_translator:av_read -> emptyreg_2:read
	wire   [31:0] emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                        // emptyreg_2:readdata -> emptyreg_2_avalon_slave_0_translator:av_readdata
	wire   [31:0] endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                     // EndTSetReg_2_avalon_slave_0_translator:av_writedata -> EndTSetReg_2:writedata
	wire    [1:0] endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address;                                       // EndTSetReg_2_avalon_slave_0_translator:av_address -> EndTSetReg_2:address
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                    // EndTSetReg_2_avalon_slave_0_translator:av_chipselect -> EndTSetReg_2:chipselect
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write;                                         // EndTSetReg_2_avalon_slave_0_translator:av_write -> EndTSetReg_2:write
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read;                                          // EndTSetReg_2_avalon_slave_0_translator:av_read -> EndTSetReg_2:read
	wire   [31:0] endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                      // EndTSetReg_2:readdata -> EndTSetReg_2_avalon_slave_0_translator:av_readdata
	wire   [31:0] fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                        // FullReg_2_avalon_slave_0_translator:av_writedata -> FullReg_2:writedata
	wire    [1:0] fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address;                                          // FullReg_2_avalon_slave_0_translator:av_address -> FullReg_2:address
	wire          fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                       // FullReg_2_avalon_slave_0_translator:av_chipselect -> FullReg_2:chipselect
	wire          fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write;                                            // FullReg_2_avalon_slave_0_translator:av_write -> FullReg_2:write
	wire          fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read;                                             // FullReg_2_avalon_slave_0_translator:av_read -> FullReg_2:read
	wire   [31:0] fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                         // FullReg_2:readdata -> FullReg_2_avalon_slave_0_translator:av_readdata
	wire   [31:0] ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                         // NTrReg_2_avalon_slave_0_translator:av_writedata -> NTrReg_2:writedata
	wire    [1:0] ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address;                                           // NTrReg_2_avalon_slave_0_translator:av_address -> NTrReg_2:address
	wire          ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                                        // NTrReg_2_avalon_slave_0_translator:av_chipselect -> NTrReg_2:chipselect
	wire          ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write;                                             // NTrReg_2_avalon_slave_0_translator:av_write -> NTrReg_2:write
	wire          ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read;                                              // NTrReg_2_avalon_slave_0_translator:av_read -> NTrReg_2:read
	wire   [31:0] ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                          // NTrReg_2:readdata -> NTrReg_2_avalon_slave_0_translator:av_readdata
	wire          dma_write_master_waitrequest;                                                                             // dma_write_master_translator:av_waitrequest -> dma:write_waitrequest
	wire   [31:0] dma_write_master_writedata;                                                                               // dma:write_writedata -> dma_write_master_translator:av_writedata
	wire   [12:0] dma_write_master_address;                                                                                 // dma:write_address -> dma_write_master_translator:av_address
	wire          dma_write_master_chipselect;                                                                              // dma:write_chipselect -> dma_write_master_translator:av_chipselect
	wire          dma_write_master_write;                                                                                   // dma:write_write_n -> dma_write_master_translator:av_write
	wire    [3:0] dma_write_master_byteenable;                                                                              // dma:write_byteenable -> dma_write_master_translator:av_byteenable
	wire          distancecore_2_avalon_master_waitrequest;                                                                 // distancecore_2_avalon_master_translator:av_waitrequest -> distancecore_2:waitrequest
	wire   [31:0] distancecore_2_avalon_master_writedata;                                                                   // distancecore_2:writedata -> distancecore_2_avalon_master_translator:av_writedata
	wire   [15:0] distancecore_2_avalon_master_address;                                                                     // distancecore_2:address -> distancecore_2_avalon_master_translator:av_address
	wire          distancecore_2_avalon_master_chipselect;                                                                  // distancecore_2:chipselect -> distancecore_2_avalon_master_translator:av_chipselect
	wire          distancecore_2_avalon_master_write;                                                                       // distancecore_2:write -> distancecore_2_avalon_master_translator:av_write
	wire          distancecore_2_avalon_master_read;                                                                        // distancecore_2:read -> distancecore_2_avalon_master_translator:av_read
	wire   [31:0] distancecore_2_avalon_master_readdata;                                                                    // distancecore_2_avalon_master_translator:av_readdata -> distancecore_2:readdata
	wire          distancecore_1_avalon_master_waitrequest;                                                                 // distancecore_1_avalon_master_translator:av_waitrequest -> distancecore_1:waitrequest
	wire   [31:0] distancecore_1_avalon_master_writedata;                                                                   // distancecore_1:writedata -> distancecore_1_avalon_master_translator:av_writedata
	wire   [15:0] distancecore_1_avalon_master_address;                                                                     // distancecore_1:address -> distancecore_1_avalon_master_translator:av_address
	wire          distancecore_1_avalon_master_chipselect;                                                                  // distancecore_1:chipselect -> distancecore_1_avalon_master_translator:av_chipselect
	wire          distancecore_1_avalon_master_write;                                                                       // distancecore_1:write -> distancecore_1_avalon_master_translator:av_write
	wire          distancecore_1_avalon_master_read;                                                                        // distancecore_1:read -> distancecore_1_avalon_master_translator:av_read
	wire   [31:0] distancecore_1_avalon_master_readdata;                                                                    // distancecore_1_avalon_master_translator:av_readdata -> distancecore_1:readdata
	wire          distancecore_0_avalon_master_waitrequest;                                                                 // distancecore_0_avalon_master_translator:av_waitrequest -> distancecore_0:waitrequest
	wire   [31:0] distancecore_0_avalon_master_writedata;                                                                   // distancecore_0:writedata -> distancecore_0_avalon_master_translator:av_writedata
	wire   [15:0] distancecore_0_avalon_master_address;                                                                     // distancecore_0:address -> distancecore_0_avalon_master_translator:av_address
	wire          distancecore_0_avalon_master_chipselect;                                                                  // distancecore_0:chipselect -> distancecore_0_avalon_master_translator:av_chipselect
	wire          distancecore_0_avalon_master_write;                                                                       // distancecore_0:write -> distancecore_0_avalon_master_translator:av_write
	wire          distancecore_0_avalon_master_read;                                                                        // distancecore_0:read -> distancecore_0_avalon_master_translator:av_read
	wire   [31:0] distancecore_0_avalon_master_readdata;                                                                    // distancecore_0_avalon_master_translator:av_readdata -> distancecore_0:readdata
	wire   [31:0] cache_0_s1_translator_avalon_anti_slave_0_writedata;                                                      // cache_0_s1_translator:av_writedata -> cache_0:writedata
	wire    [8:0] cache_0_s1_translator_avalon_anti_slave_0_address;                                                        // cache_0_s1_translator:av_address -> cache_0:address
	wire          cache_0_s1_translator_avalon_anti_slave_0_chipselect;                                                     // cache_0_s1_translator:av_chipselect -> cache_0:chipselect
	wire          cache_0_s1_translator_avalon_anti_slave_0_clken;                                                          // cache_0_s1_translator:av_clken -> cache_0:clken
	wire          cache_0_s1_translator_avalon_anti_slave_0_write;                                                          // cache_0_s1_translator:av_write -> cache_0:write
	wire   [31:0] cache_0_s1_translator_avalon_anti_slave_0_readdata;                                                       // cache_0:readdata -> cache_0_s1_translator:av_readdata
	wire    [3:0] cache_0_s1_translator_avalon_anti_slave_0_byteenable;                                                     // cache_0_s1_translator:av_byteenable -> cache_0:byteenable
	wire   [31:0] cache_1_s1_translator_avalon_anti_slave_0_writedata;                                                      // cache_1_s1_translator:av_writedata -> cache_1:writedata
	wire    [8:0] cache_1_s1_translator_avalon_anti_slave_0_address;                                                        // cache_1_s1_translator:av_address -> cache_1:address
	wire          cache_1_s1_translator_avalon_anti_slave_0_chipselect;                                                     // cache_1_s1_translator:av_chipselect -> cache_1:chipselect
	wire          cache_1_s1_translator_avalon_anti_slave_0_clken;                                                          // cache_1_s1_translator:av_clken -> cache_1:clken
	wire          cache_1_s1_translator_avalon_anti_slave_0_write;                                                          // cache_1_s1_translator:av_write -> cache_1:write
	wire   [31:0] cache_1_s1_translator_avalon_anti_slave_0_readdata;                                                       // cache_1:readdata -> cache_1_s1_translator:av_readdata
	wire    [3:0] cache_1_s1_translator_avalon_anti_slave_0_byteenable;                                                     // cache_1_s1_translator:av_byteenable -> cache_1:byteenable
	wire   [31:0] cache_2_s1_translator_avalon_anti_slave_0_writedata;                                                      // cache_2_s1_translator:av_writedata -> cache_2:writedata
	wire    [8:0] cache_2_s1_translator_avalon_anti_slave_0_address;                                                        // cache_2_s1_translator:av_address -> cache_2:address
	wire          cache_2_s1_translator_avalon_anti_slave_0_chipselect;                                                     // cache_2_s1_translator:av_chipselect -> cache_2:chipselect
	wire          cache_2_s1_translator_avalon_anti_slave_0_clken;                                                          // cache_2_s1_translator:av_clken -> cache_2:clken
	wire          cache_2_s1_translator_avalon_anti_slave_0_write;                                                          // cache_2_s1_translator:av_write -> cache_2:write
	wire   [31:0] cache_2_s1_translator_avalon_anti_slave_0_readdata;                                                       // cache_2:readdata -> cache_2_s1_translator:av_readdata
	wire    [3:0] cache_2_s1_translator_avalon_anti_slave_0_byteenable;                                                     // cache_2_s1_translator:av_byteenable -> cache_2:byteenable
	wire          distancecore_0_avalon_master_1_waitrequest;                                                               // distancecore_0_avalon_master_1_translator:av_waitrequest -> distancecore_0:waitrequest1
	wire   [31:0] distancecore_0_avalon_master_1_writedata;                                                                 // distancecore_0:writedata1 -> distancecore_0_avalon_master_1_translator:av_writedata
	wire   [15:0] distancecore_0_avalon_master_1_address;                                                                   // distancecore_0:address1 -> distancecore_0_avalon_master_1_translator:av_address
	wire          distancecore_0_avalon_master_1_chipselect;                                                                // distancecore_0:chipselect1 -> distancecore_0_avalon_master_1_translator:av_chipselect
	wire          distancecore_0_avalon_master_1_write;                                                                     // distancecore_0:write1 -> distancecore_0_avalon_master_1_translator:av_write
	wire          distancecore_0_avalon_master_1_read;                                                                      // distancecore_0:read1 -> distancecore_0_avalon_master_1_translator:av_read
	wire   [31:0] distancecore_0_avalon_master_1_readdata;                                                                  // distancecore_0_avalon_master_1_translator:av_readdata -> distancecore_0:readdata1
	wire   [31:0] cache_0_s2_translator_avalon_anti_slave_0_writedata;                                                      // cache_0_s2_translator:av_writedata -> cache_0:writedata2
	wire    [8:0] cache_0_s2_translator_avalon_anti_slave_0_address;                                                        // cache_0_s2_translator:av_address -> cache_0:address2
	wire          cache_0_s2_translator_avalon_anti_slave_0_chipselect;                                                     // cache_0_s2_translator:av_chipselect -> cache_0:chipselect2
	wire          cache_0_s2_translator_avalon_anti_slave_0_clken;                                                          // cache_0_s2_translator:av_clken -> cache_0:clken2
	wire          cache_0_s2_translator_avalon_anti_slave_0_write;                                                          // cache_0_s2_translator:av_write -> cache_0:write2
	wire   [31:0] cache_0_s2_translator_avalon_anti_slave_0_readdata;                                                       // cache_0:readdata2 -> cache_0_s2_translator:av_readdata
	wire    [3:0] cache_0_s2_translator_avalon_anti_slave_0_byteenable;                                                     // cache_0_s2_translator:av_byteenable -> cache_0:byteenable2
	wire          distancecore_1_avalon_master_1_waitrequest;                                                               // distancecore_1_avalon_master_1_translator:av_waitrequest -> distancecore_1:waitrequest1
	wire   [31:0] distancecore_1_avalon_master_1_writedata;                                                                 // distancecore_1:writedata1 -> distancecore_1_avalon_master_1_translator:av_writedata
	wire   [15:0] distancecore_1_avalon_master_1_address;                                                                   // distancecore_1:address1 -> distancecore_1_avalon_master_1_translator:av_address
	wire          distancecore_1_avalon_master_1_chipselect;                                                                // distancecore_1:chipselect1 -> distancecore_1_avalon_master_1_translator:av_chipselect
	wire          distancecore_1_avalon_master_1_write;                                                                     // distancecore_1:write1 -> distancecore_1_avalon_master_1_translator:av_write
	wire          distancecore_1_avalon_master_1_read;                                                                      // distancecore_1:read1 -> distancecore_1_avalon_master_1_translator:av_read
	wire   [31:0] distancecore_1_avalon_master_1_readdata;                                                                  // distancecore_1_avalon_master_1_translator:av_readdata -> distancecore_1:readdata1
	wire   [31:0] cache_1_s2_translator_avalon_anti_slave_0_writedata;                                                      // cache_1_s2_translator:av_writedata -> cache_1:writedata2
	wire    [8:0] cache_1_s2_translator_avalon_anti_slave_0_address;                                                        // cache_1_s2_translator:av_address -> cache_1:address2
	wire          cache_1_s2_translator_avalon_anti_slave_0_chipselect;                                                     // cache_1_s2_translator:av_chipselect -> cache_1:chipselect2
	wire          cache_1_s2_translator_avalon_anti_slave_0_clken;                                                          // cache_1_s2_translator:av_clken -> cache_1:clken2
	wire          cache_1_s2_translator_avalon_anti_slave_0_write;                                                          // cache_1_s2_translator:av_write -> cache_1:write2
	wire   [31:0] cache_1_s2_translator_avalon_anti_slave_0_readdata;                                                       // cache_1:readdata2 -> cache_1_s2_translator:av_readdata
	wire    [3:0] cache_1_s2_translator_avalon_anti_slave_0_byteenable;                                                     // cache_1_s2_translator:av_byteenable -> cache_1:byteenable2
	wire          distancecore_2_avalon_master_1_waitrequest;                                                               // distancecore_2_avalon_master_1_translator:av_waitrequest -> distancecore_2:waitrequest1
	wire   [31:0] distancecore_2_avalon_master_1_writedata;                                                                 // distancecore_2:writedata1 -> distancecore_2_avalon_master_1_translator:av_writedata
	wire   [15:0] distancecore_2_avalon_master_1_address;                                                                   // distancecore_2:address1 -> distancecore_2_avalon_master_1_translator:av_address
	wire          distancecore_2_avalon_master_1_chipselect;                                                                // distancecore_2:chipselect1 -> distancecore_2_avalon_master_1_translator:av_chipselect
	wire          distancecore_2_avalon_master_1_write;                                                                     // distancecore_2:write1 -> distancecore_2_avalon_master_1_translator:av_write
	wire          distancecore_2_avalon_master_1_read;                                                                      // distancecore_2:read1 -> distancecore_2_avalon_master_1_translator:av_read
	wire   [31:0] distancecore_2_avalon_master_1_readdata;                                                                  // distancecore_2_avalon_master_1_translator:av_readdata -> distancecore_2:readdata1
	wire   [31:0] cache_2_s2_translator_avalon_anti_slave_0_writedata;                                                      // cache_2_s2_translator:av_writedata -> cache_2:writedata2
	wire    [8:0] cache_2_s2_translator_avalon_anti_slave_0_address;                                                        // cache_2_s2_translator:av_address -> cache_2:address2
	wire          cache_2_s2_translator_avalon_anti_slave_0_chipselect;                                                     // cache_2_s2_translator:av_chipselect -> cache_2:chipselect2
	wire          cache_2_s2_translator_avalon_anti_slave_0_clken;                                                          // cache_2_s2_translator:av_clken -> cache_2:clken2
	wire          cache_2_s2_translator_avalon_anti_slave_0_write;                                                          // cache_2_s2_translator:av_write -> cache_2:write2
	wire   [31:0] cache_2_s2_translator_avalon_anti_slave_0_readdata;                                                       // cache_2:readdata2 -> cache_2_s2_translator:av_readdata
	wire    [3:0] cache_2_s2_translator_avalon_anti_slave_0_byteenable;                                                     // cache_2_s2_translator:av_byteenable -> cache_2:byteenable2
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                                // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount;                                 // cpu_0_instruction_master_translator:uav_burstcount -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_writedata;                                  // cpu_0_instruction_master_translator:uav_writedata -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] cpu_0_instruction_master_translator_avalon_universal_master_0_address;                                    // cpu_0_instruction_master_translator:uav_address -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_lock;                                       // cpu_0_instruction_master_translator:uav_lock -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_write;                                      // cpu_0_instruction_master_translator:uav_write -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_read;                                       // cpu_0_instruction_master_translator:uav_read -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_0_instruction_master_translator_avalon_universal_master_0_readdata;                                   // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_instruction_master_translator:uav_readdata
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                                // cpu_0_instruction_master_translator:uav_debugaccess -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable;                                 // cpu_0_instruction_master_translator:uav_byteenable -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_instruction_master_translator:uav_readdatavalid
	wire          cpu_0_data_master_translator_avalon_universal_master_0_waitrequest;                                       // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_0_data_master_translator_avalon_universal_master_0_burstcount;                                        // cpu_0_data_master_translator:uav_burstcount -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_0_data_master_translator_avalon_universal_master_0_writedata;                                         // cpu_0_data_master_translator:uav_writedata -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] cpu_0_data_master_translator_avalon_universal_master_0_address;                                           // cpu_0_data_master_translator:uav_address -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_0_data_master_translator_avalon_universal_master_0_lock;                                              // cpu_0_data_master_translator:uav_lock -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_0_data_master_translator_avalon_universal_master_0_write;                                             // cpu_0_data_master_translator:uav_write -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_0_data_master_translator_avalon_universal_master_0_read;                                              // cpu_0_data_master_translator:uav_read -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_0_data_master_translator_avalon_universal_master_0_readdata;                                          // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_data_master_translator:uav_readdata
	wire          cpu_0_data_master_translator_avalon_universal_master_0_debugaccess;                                       // cpu_0_data_master_translator:uav_debugaccess -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_0_data_master_translator_avalon_universal_master_0_byteenable;                                        // cpu_0_data_master_translator:uav_byteenable -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                     // cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_data_master_translator:uav_readdatavalid
	wire          dma_read_master_translator_avalon_universal_master_0_waitrequest;                                         // dma_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_read_master_translator:uav_waitrequest
	wire    [2:0] dma_read_master_translator_avalon_universal_master_0_burstcount;                                          // dma_read_master_translator:uav_burstcount -> dma_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_read_master_translator_avalon_universal_master_0_writedata;                                           // dma_read_master_translator:uav_writedata -> dma_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [25:0] dma_read_master_translator_avalon_universal_master_0_address;                                             // dma_read_master_translator:uav_address -> dma_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_read_master_translator_avalon_universal_master_0_lock;                                                // dma_read_master_translator:uav_lock -> dma_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_read_master_translator_avalon_universal_master_0_write;                                               // dma_read_master_translator:uav_write -> dma_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_read_master_translator_avalon_universal_master_0_read;                                                // dma_read_master_translator:uav_read -> dma_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_read_master_translator_avalon_universal_master_0_readdata;                                            // dma_read_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_read_master_translator:uav_readdata
	wire          dma_read_master_translator_avalon_universal_master_0_debugaccess;                                         // dma_read_master_translator:uav_debugaccess -> dma_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_read_master_translator_avalon_universal_master_0_byteenable;                                          // dma_read_master_translator:uav_byteenable -> dma_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_read_master_translator_avalon_universal_master_0_readdatavalid;                                       // dma_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_read_master_translator:uav_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire   [25:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // dma_control_port_slave_translator:uav_waitrequest -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dma_control_port_slave_translator:uav_burstcount
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                            // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dma_control_port_slave_translator:uav_writedata
	wire   [25:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                              // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> dma_control_port_slave_translator:uav_address
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                                // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> dma_control_port_slave_translator:uav_write
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> dma_control_port_slave_translator:uav_lock
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> dma_control_port_slave_translator:uav_read
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                             // dma_control_port_slave_translator:uav_readdata -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // dma_control_port_slave_translator:uav_readdatavalid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dma_control_port_slave_translator:uav_debugaccess
	wire    [3:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // dma_control_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dma_control_port_slave_translator:uav_byteenable
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                          // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [25:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // pio_0_s1_translator:uav_waitrequest -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_0_s1_translator:uav_burstcount
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_0_s1_translator:uav_writedata
	wire   [25:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                            // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_0_s1_translator:uav_address
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                              // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_0_s1_translator:uav_write
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                               // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_0_s1_translator:uav_lock
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                               // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_0_s1_translator:uav_read
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // pio_0_s1_translator:uav_readdata -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // pio_0_s1_translator:uav_readdatavalid -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_0_s1_translator:uav_debugaccess
	wire    [3:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_0_s1_translator:uav_byteenable
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // usbFIFOCtrl_0_avalon_slave_0_translator:uav_waitrequest -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> usbFIFOCtrl_0_avalon_slave_0_translator:uav_burstcount
	wire   [15:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                      // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> usbFIFOCtrl_0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                        // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> usbFIFOCtrl_0_avalon_slave_0_translator:uav_address
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                          // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> usbFIFOCtrl_0_avalon_slave_0_translator:uav_write
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                           // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> usbFIFOCtrl_0_avalon_slave_0_translator:uav_lock
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                           // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> usbFIFOCtrl_0_avalon_slave_0_translator:uav_read
	wire   [15:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                       // usbFIFOCtrl_0_avalon_slave_0_translator:uav_readdata -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // usbFIFOCtrl_0_avalon_slave_0_translator:uav_readdatavalid -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> usbFIFOCtrl_0_avalon_slave_0_translator:uav_debugaccess
	wire    [1:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> usbFIFOCtrl_0_avalon_slave_0_translator:uav_byteenable
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                    // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [15:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;              // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [15:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;               // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;              // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // sdram_controller_s1_translator:uav_waitrequest -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_controller_s1_translator:uav_burstcount
	wire   [31:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_controller_s1_translator:uav_writedata
	wire   [25:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_controller_s1_translator:uav_address
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_controller_s1_translator:uav_write
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_controller_s1_translator:uav_lock
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_controller_s1_translator:uav_read
	wire   [31:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // sdram_controller_s1_translator:uav_readdata -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // sdram_controller_s1_translator:uav_readdatavalid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_controller_s1_translator:uav_debugaccess
	wire    [3:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // sdram_controller_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_controller_s1_translator:uav_byteenable
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // performance_counter_0_control_slave_translator:uav_waitrequest -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_0_control_slave_translator:uav_burstcount
	wire   [31:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_0_control_slave_translator:uav_writedata
	wire   [25:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_0_control_slave_translator:uav_address
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_0_control_slave_translator:uav_write
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_0_control_slave_translator:uav_lock
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_0_control_slave_translator:uav_read
	wire   [31:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // performance_counter_0_control_slave_translator:uav_readdata -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // performance_counter_0_control_slave_translator:uav_readdatavalid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_0_control_slave_translator:uav_debugaccess
	wire    [3:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_0_control_slave_translator:uav_byteenable
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // NDimReg_avalon_slave_0_translator:uav_waitrequest -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> NDimReg_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                            // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> NDimReg_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                              // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> NDimReg_avalon_slave_0_translator:uav_address
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> NDimReg_avalon_slave_0_translator:uav_write
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                 // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> NDimReg_avalon_slave_0_translator:uav_lock
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                 // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> NDimReg_avalon_slave_0_translator:uav_read
	wire   [31:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                             // NDimReg_avalon_slave_0_translator:uav_readdata -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // NDimReg_avalon_slave_0_translator:uav_readdatavalid -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NDimReg_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> NDimReg_avalon_slave_0_translator:uav_byteenable
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                          // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                    // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                     // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                    // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // EndTSetReg_0_avalon_slave_0_translator:uav_waitrequest -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> EndTSetReg_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                       // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> EndTSetReg_0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                         // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> EndTSetReg_0_avalon_slave_0_translator:uav_address
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                           // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> EndTSetReg_0_avalon_slave_0_translator:uav_write
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                            // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> EndTSetReg_0_avalon_slave_0_translator:uav_lock
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                            // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> EndTSetReg_0_avalon_slave_0_translator:uav_read
	wire   [31:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                        // EndTSetReg_0_avalon_slave_0_translator:uav_readdata -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // EndTSetReg_0_avalon_slave_0_translator:uav_readdatavalid -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> EndTSetReg_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> EndTSetReg_0_avalon_slave_0_translator:uav_byteenable
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                     // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;               // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;               // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // FullReg_0_avalon_slave_0_translator:uav_waitrequest -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> FullReg_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                          // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> FullReg_0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                            // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> FullReg_0_avalon_slave_0_translator:uav_address
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                              // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> FullReg_0_avalon_slave_0_translator:uav_write
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                               // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> FullReg_0_avalon_slave_0_translator:uav_lock
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                               // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> FullReg_0_avalon_slave_0_translator:uav_read
	wire   [31:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                           // FullReg_0_avalon_slave_0_translator:uav_readdata -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // FullReg_0_avalon_slave_0_translator:uav_readdatavalid -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FullReg_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> FullReg_0_avalon_slave_0_translator:uav_byteenable
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                        // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // FullReg_1_avalon_slave_0_translator:uav_waitrequest -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> FullReg_1_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                          // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> FullReg_1_avalon_slave_0_translator:uav_writedata
	wire   [25:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                            // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> FullReg_1_avalon_slave_0_translator:uav_address
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                              // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> FullReg_1_avalon_slave_0_translator:uav_write
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                               // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> FullReg_1_avalon_slave_0_translator:uav_lock
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                               // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> FullReg_1_avalon_slave_0_translator:uav_read
	wire   [31:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                           // FullReg_1_avalon_slave_0_translator:uav_readdata -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // FullReg_1_avalon_slave_0_translator:uav_readdatavalid -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FullReg_1_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> FullReg_1_avalon_slave_0_translator:uav_byteenable
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                        // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // NTrReg_0_avalon_slave_0_translator:uav_waitrequest -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> NTrReg_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                           // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> NTrReg_0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                             // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> NTrReg_0_avalon_slave_0_translator:uav_address
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                               // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> NTrReg_0_avalon_slave_0_translator:uav_write
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> NTrReg_0_avalon_slave_0_translator:uav_lock
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> NTrReg_0_avalon_slave_0_translator:uav_read
	wire   [31:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                            // NTrReg_0_avalon_slave_0_translator:uav_readdata -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // NTrReg_0_avalon_slave_0_translator:uav_readdatavalid -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NTrReg_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> NTrReg_0_avalon_slave_0_translator:uav_byteenable
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                         // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                   // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                    // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                   // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // NTrReg_1_avalon_slave_0_translator:uav_waitrequest -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> NTrReg_1_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                           // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> NTrReg_1_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                             // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> NTrReg_1_avalon_slave_0_translator:uav_address
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                               // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> NTrReg_1_avalon_slave_0_translator:uav_write
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> NTrReg_1_avalon_slave_0_translator:uav_lock
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> NTrReg_1_avalon_slave_0_translator:uav_read
	wire   [31:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                            // NTrReg_1_avalon_slave_0_translator:uav_readdata -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // NTrReg_1_avalon_slave_0_translator:uav_readdatavalid -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NTrReg_1_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> NTrReg_1_avalon_slave_0_translator:uav_byteenable
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                         // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                   // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                    // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                   // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // emptyreg_0_avalon_slave_0_translator:uav_waitrequest -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> emptyreg_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                         // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> emptyreg_0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                           // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> emptyreg_0_avalon_slave_0_translator:uav_address
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                             // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> emptyreg_0_avalon_slave_0_translator:uav_write
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                              // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> emptyreg_0_avalon_slave_0_translator:uav_lock
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                              // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> emptyreg_0_avalon_slave_0_translator:uav_read
	wire   [31:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                          // emptyreg_0_avalon_slave_0_translator:uav_readdata -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // emptyreg_0_avalon_slave_0_translator:uav_readdatavalid -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> emptyreg_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> emptyreg_0_avalon_slave_0_translator:uav_byteenable
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                       // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // emptyreg_1_avalon_slave_0_translator:uav_waitrequest -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> emptyreg_1_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                         // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> emptyreg_1_avalon_slave_0_translator:uav_writedata
	wire   [25:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                           // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> emptyreg_1_avalon_slave_0_translator:uav_address
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                             // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> emptyreg_1_avalon_slave_0_translator:uav_write
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                              // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> emptyreg_1_avalon_slave_0_translator:uav_lock
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                              // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> emptyreg_1_avalon_slave_0_translator:uav_read
	wire   [31:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                          // emptyreg_1_avalon_slave_0_translator:uav_readdata -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // emptyreg_1_avalon_slave_0_translator:uav_readdatavalid -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> emptyreg_1_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> emptyreg_1_avalon_slave_0_translator:uav_byteenable
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                       // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // EndTSetReg_1_avalon_slave_0_translator:uav_waitrequest -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> EndTSetReg_1_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                       // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> EndTSetReg_1_avalon_slave_0_translator:uav_writedata
	wire   [25:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                         // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> EndTSetReg_1_avalon_slave_0_translator:uav_address
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                           // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> EndTSetReg_1_avalon_slave_0_translator:uav_write
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                            // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> EndTSetReg_1_avalon_slave_0_translator:uav_lock
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                            // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> EndTSetReg_1_avalon_slave_0_translator:uav_read
	wire   [31:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                        // EndTSetReg_1_avalon_slave_0_translator:uav_readdata -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // EndTSetReg_1_avalon_slave_0_translator:uav_readdatavalid -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> EndTSetReg_1_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> EndTSetReg_1_avalon_slave_0_translator:uav_byteenable
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                     // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;               // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;               // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // baseqaddr_0_avalon_slave_0_translator:uav_waitrequest -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> baseqaddr_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                        // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> baseqaddr_0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                          // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> baseqaddr_0_avalon_slave_0_translator:uav_address
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                            // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> baseqaddr_0_avalon_slave_0_translator:uav_write
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                             // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> baseqaddr_0_avalon_slave_0_translator:uav_lock
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                             // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> baseqaddr_0_avalon_slave_0_translator:uav_read
	wire   [31:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                         // baseqaddr_0_avalon_slave_0_translator:uav_readdata -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // baseqaddr_0_avalon_slave_0_translator:uav_readdatavalid -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> baseqaddr_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> baseqaddr_0_avalon_slave_0_translator:uav_byteenable
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                      // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // skipaddrreg_0_avalon_slave_0_translator:uav_waitrequest -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> skipaddrreg_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                      // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> skipaddrreg_0_avalon_slave_0_translator:uav_writedata
	wire   [25:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                        // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> skipaddrreg_0_avalon_slave_0_translator:uav_address
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                          // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> skipaddrreg_0_avalon_slave_0_translator:uav_write
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                           // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> skipaddrreg_0_avalon_slave_0_translator:uav_lock
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                           // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> skipaddrreg_0_avalon_slave_0_translator:uav_read
	wire   [31:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                       // skipaddrreg_0_avalon_slave_0_translator:uav_readdata -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // skipaddrreg_0_avalon_slave_0_translator:uav_readdatavalid -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> skipaddrreg_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> skipaddrreg_0_avalon_slave_0_translator:uav_byteenable
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                    // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;              // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;               // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;              // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // knnclasscore_avalon_slave_0_translator:uav_waitrequest -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> knnclasscore_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                       // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> knnclasscore_avalon_slave_0_translator:uav_writedata
	wire   [25:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                         // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> knnclasscore_avalon_slave_0_translator:uav_address
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                           // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> knnclasscore_avalon_slave_0_translator:uav_write
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                            // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> knnclasscore_avalon_slave_0_translator:uav_lock
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                            // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> knnclasscore_avalon_slave_0_translator:uav_read
	wire   [31:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                        // knnclasscore_avalon_slave_0_translator:uav_readdata -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // knnclasscore_avalon_slave_0_translator:uav_readdatavalid -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> knnclasscore_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> knnclasscore_avalon_slave_0_translator:uav_byteenable
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                     // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;               // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;               // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // emptyreg_2_avalon_slave_0_translator:uav_waitrequest -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> emptyreg_2_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                         // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> emptyreg_2_avalon_slave_0_translator:uav_writedata
	wire   [25:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                           // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> emptyreg_2_avalon_slave_0_translator:uav_address
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                             // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> emptyreg_2_avalon_slave_0_translator:uav_write
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                              // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> emptyreg_2_avalon_slave_0_translator:uav_lock
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                              // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> emptyreg_2_avalon_slave_0_translator:uav_read
	wire   [31:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                          // emptyreg_2_avalon_slave_0_translator:uav_readdata -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // emptyreg_2_avalon_slave_0_translator:uav_readdatavalid -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> emptyreg_2_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> emptyreg_2_avalon_slave_0_translator:uav_byteenable
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                       // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                 // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                  // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                 // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // EndTSetReg_2_avalon_slave_0_translator:uav_waitrequest -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> EndTSetReg_2_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                       // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> EndTSetReg_2_avalon_slave_0_translator:uav_writedata
	wire   [25:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                         // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> EndTSetReg_2_avalon_slave_0_translator:uav_address
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                           // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> EndTSetReg_2_avalon_slave_0_translator:uav_write
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                            // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> EndTSetReg_2_avalon_slave_0_translator:uav_lock
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                            // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> EndTSetReg_2_avalon_slave_0_translator:uav_read
	wire   [31:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                        // EndTSetReg_2_avalon_slave_0_translator:uav_readdata -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // EndTSetReg_2_avalon_slave_0_translator:uav_readdatavalid -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> EndTSetReg_2_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> EndTSetReg_2_avalon_slave_0_translator:uav_byteenable
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                     // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;               // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;               // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // FullReg_2_avalon_slave_0_translator:uav_waitrequest -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> FullReg_2_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                          // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> FullReg_2_avalon_slave_0_translator:uav_writedata
	wire   [25:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                            // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> FullReg_2_avalon_slave_0_translator:uav_address
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                              // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> FullReg_2_avalon_slave_0_translator:uav_write
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                               // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> FullReg_2_avalon_slave_0_translator:uav_lock
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                               // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> FullReg_2_avalon_slave_0_translator:uav_read
	wire   [31:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                           // FullReg_2_avalon_slave_0_translator:uav_readdata -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // FullReg_2_avalon_slave_0_translator:uav_readdatavalid -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> FullReg_2_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> FullReg_2_avalon_slave_0_translator:uav_byteenable
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                        // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                  // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                   // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                  // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // NTrReg_2_avalon_slave_0_translator:uav_waitrequest -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> NTrReg_2_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                           // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> NTrReg_2_avalon_slave_0_translator:uav_writedata
	wire   [25:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                             // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> NTrReg_2_avalon_slave_0_translator:uav_address
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                               // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> NTrReg_2_avalon_slave_0_translator:uav_write
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> NTrReg_2_avalon_slave_0_translator:uav_lock
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> NTrReg_2_avalon_slave_0_translator:uav_read
	wire   [31:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                            // NTrReg_2_avalon_slave_0_translator:uav_readdata -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // NTrReg_2_avalon_slave_0_translator:uav_readdatavalid -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NTrReg_2_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> NTrReg_2_avalon_slave_0_translator:uav_byteenable
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [103:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                         // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [103:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                   // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                    // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                   // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dma_write_master_translator_avalon_universal_master_0_waitrequest;                                        // dma_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_write_master_translator:uav_waitrequest
	wire    [2:0] dma_write_master_translator_avalon_universal_master_0_burstcount;                                         // dma_write_master_translator:uav_burstcount -> dma_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] dma_write_master_translator_avalon_universal_master_0_writedata;                                          // dma_write_master_translator:uav_writedata -> dma_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] dma_write_master_translator_avalon_universal_master_0_address;                                            // dma_write_master_translator:uav_address -> dma_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_write_master_translator_avalon_universal_master_0_lock;                                               // dma_write_master_translator:uav_lock -> dma_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_write_master_translator_avalon_universal_master_0_write;                                              // dma_write_master_translator:uav_write -> dma_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_write_master_translator_avalon_universal_master_0_read;                                               // dma_write_master_translator:uav_read -> dma_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] dma_write_master_translator_avalon_universal_master_0_readdata;                                           // dma_write_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_write_master_translator:uav_readdata
	wire          dma_write_master_translator_avalon_universal_master_0_debugaccess;                                        // dma_write_master_translator:uav_debugaccess -> dma_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] dma_write_master_translator_avalon_universal_master_0_byteenable;                                         // dma_write_master_translator:uav_byteenable -> dma_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_write_master_translator_avalon_universal_master_0_readdatavalid;                                      // dma_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_write_master_translator:uav_readdatavalid
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_waitrequest;                            // distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> distancecore_2_avalon_master_translator:uav_waitrequest
	wire    [2:0] distancecore_2_avalon_master_translator_avalon_universal_master_0_burstcount;                             // distancecore_2_avalon_master_translator:uav_burstcount -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] distancecore_2_avalon_master_translator_avalon_universal_master_0_writedata;                              // distancecore_2_avalon_master_translator:uav_writedata -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] distancecore_2_avalon_master_translator_avalon_universal_master_0_address;                                // distancecore_2_avalon_master_translator:uav_address -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_lock;                                   // distancecore_2_avalon_master_translator:uav_lock -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_write;                                  // distancecore_2_avalon_master_translator:uav_write -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_read;                                   // distancecore_2_avalon_master_translator:uav_read -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] distancecore_2_avalon_master_translator_avalon_universal_master_0_readdata;                               // distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> distancecore_2_avalon_master_translator:uav_readdata
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_debugaccess;                            // distancecore_2_avalon_master_translator:uav_debugaccess -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] distancecore_2_avalon_master_translator_avalon_universal_master_0_byteenable;                             // distancecore_2_avalon_master_translator:uav_byteenable -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_readdatavalid;                          // distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> distancecore_2_avalon_master_translator:uav_readdatavalid
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_waitrequest;                            // distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> distancecore_1_avalon_master_translator:uav_waitrequest
	wire    [2:0] distancecore_1_avalon_master_translator_avalon_universal_master_0_burstcount;                             // distancecore_1_avalon_master_translator:uav_burstcount -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] distancecore_1_avalon_master_translator_avalon_universal_master_0_writedata;                              // distancecore_1_avalon_master_translator:uav_writedata -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] distancecore_1_avalon_master_translator_avalon_universal_master_0_address;                                // distancecore_1_avalon_master_translator:uav_address -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_lock;                                   // distancecore_1_avalon_master_translator:uav_lock -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_write;                                  // distancecore_1_avalon_master_translator:uav_write -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_read;                                   // distancecore_1_avalon_master_translator:uav_read -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] distancecore_1_avalon_master_translator_avalon_universal_master_0_readdata;                               // distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> distancecore_1_avalon_master_translator:uav_readdata
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_debugaccess;                            // distancecore_1_avalon_master_translator:uav_debugaccess -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] distancecore_1_avalon_master_translator_avalon_universal_master_0_byteenable;                             // distancecore_1_avalon_master_translator:uav_byteenable -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_readdatavalid;                          // distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> distancecore_1_avalon_master_translator:uav_readdatavalid
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_waitrequest;                            // distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> distancecore_0_avalon_master_translator:uav_waitrequest
	wire    [2:0] distancecore_0_avalon_master_translator_avalon_universal_master_0_burstcount;                             // distancecore_0_avalon_master_translator:uav_burstcount -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] distancecore_0_avalon_master_translator_avalon_universal_master_0_writedata;                              // distancecore_0_avalon_master_translator:uav_writedata -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] distancecore_0_avalon_master_translator_avalon_universal_master_0_address;                                // distancecore_0_avalon_master_translator:uav_address -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_lock;                                   // distancecore_0_avalon_master_translator:uav_lock -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_write;                                  // distancecore_0_avalon_master_translator:uav_write -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_read;                                   // distancecore_0_avalon_master_translator:uav_read -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] distancecore_0_avalon_master_translator_avalon_universal_master_0_readdata;                               // distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> distancecore_0_avalon_master_translator:uav_readdata
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_debugaccess;                            // distancecore_0_avalon_master_translator:uav_debugaccess -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] distancecore_0_avalon_master_translator_avalon_universal_master_0_byteenable;                             // distancecore_0_avalon_master_translator:uav_byteenable -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_readdatavalid;                          // distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> distancecore_0_avalon_master_translator:uav_readdatavalid
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // cache_0_s1_translator:uav_waitrequest -> cache_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cache_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // cache_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> cache_0_s1_translator:uav_burstcount
	wire   [31:0] cache_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // cache_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> cache_0_s1_translator:uav_writedata
	wire   [15:0] cache_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // cache_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> cache_0_s1_translator:uav_address
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // cache_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> cache_0_s1_translator:uav_write
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // cache_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> cache_0_s1_translator:uav_lock
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // cache_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> cache_0_s1_translator:uav_read
	wire   [31:0] cache_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // cache_0_s1_translator:uav_readdata -> cache_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // cache_0_s1_translator:uav_readdatavalid -> cache_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // cache_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cache_0_s1_translator:uav_debugaccess
	wire    [3:0] cache_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // cache_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> cache_0_s1_translator:uav_byteenable
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // cache_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // cache_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // cache_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [87:0] cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // cache_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cache_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cache_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cache_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cache_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [87:0] cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cache_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // cache_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // cache_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // cache_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cache_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cache_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cache_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // cache_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // cache_1_s1_translator:uav_waitrequest -> cache_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cache_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // cache_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> cache_1_s1_translator:uav_burstcount
	wire   [31:0] cache_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // cache_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> cache_1_s1_translator:uav_writedata
	wire   [15:0] cache_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // cache_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> cache_1_s1_translator:uav_address
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // cache_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> cache_1_s1_translator:uav_write
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // cache_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> cache_1_s1_translator:uav_lock
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // cache_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> cache_1_s1_translator:uav_read
	wire   [31:0] cache_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // cache_1_s1_translator:uav_readdata -> cache_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // cache_1_s1_translator:uav_readdatavalid -> cache_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // cache_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cache_1_s1_translator:uav_debugaccess
	wire    [3:0] cache_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // cache_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> cache_1_s1_translator:uav_byteenable
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // cache_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // cache_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // cache_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [87:0] cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // cache_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cache_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cache_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cache_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cache_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [87:0] cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cache_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // cache_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // cache_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // cache_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cache_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cache_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cache_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // cache_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // cache_2_s1_translator:uav_waitrequest -> cache_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cache_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // cache_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> cache_2_s1_translator:uav_burstcount
	wire   [31:0] cache_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // cache_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> cache_2_s1_translator:uav_writedata
	wire   [15:0] cache_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                          // cache_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> cache_2_s1_translator:uav_address
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                            // cache_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> cache_2_s1_translator:uav_write
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                             // cache_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> cache_2_s1_translator:uav_lock
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                             // cache_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> cache_2_s1_translator:uav_read
	wire   [31:0] cache_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // cache_2_s1_translator:uav_readdata -> cache_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // cache_2_s1_translator:uav_readdatavalid -> cache_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // cache_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cache_2_s1_translator:uav_debugaccess
	wire    [3:0] cache_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // cache_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> cache_2_s1_translator:uav_byteenable
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // cache_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // cache_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // cache_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [87:0] cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // cache_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cache_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cache_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cache_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cache_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [87:0] cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cache_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // cache_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // cache_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // cache_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cache_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cache_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cache_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // cache_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_waitrequest;                          // distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_waitrequest -> distancecore_0_avalon_master_1_translator:uav_waitrequest
	wire    [2:0] distancecore_0_avalon_master_1_translator_avalon_universal_master_0_burstcount;                           // distancecore_0_avalon_master_1_translator:uav_burstcount -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] distancecore_0_avalon_master_1_translator_avalon_universal_master_0_writedata;                            // distancecore_0_avalon_master_1_translator:uav_writedata -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] distancecore_0_avalon_master_1_translator_avalon_universal_master_0_address;                              // distancecore_0_avalon_master_1_translator:uav_address -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_address
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_lock;                                 // distancecore_0_avalon_master_1_translator:uav_lock -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_lock
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_write;                                // distancecore_0_avalon_master_1_translator:uav_write -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_write
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_read;                                 // distancecore_0_avalon_master_1_translator:uav_read -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] distancecore_0_avalon_master_1_translator_avalon_universal_master_0_readdata;                             // distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_readdata -> distancecore_0_avalon_master_1_translator:uav_readdata
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_debugaccess;                          // distancecore_0_avalon_master_1_translator:uav_debugaccess -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] distancecore_0_avalon_master_1_translator_avalon_universal_master_0_byteenable;                           // distancecore_0_avalon_master_1_translator:uav_byteenable -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_byteenable
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_readdatavalid;                        // distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:av_readdatavalid -> distancecore_0_avalon_master_1_translator:uav_readdatavalid
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // cache_0_s2_translator:uav_waitrequest -> cache_0_s2_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cache_0_s2_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // cache_0_s2_translator_avalon_universal_slave_0_agent:m0_burstcount -> cache_0_s2_translator:uav_burstcount
	wire   [31:0] cache_0_s2_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // cache_0_s2_translator_avalon_universal_slave_0_agent:m0_writedata -> cache_0_s2_translator:uav_writedata
	wire   [15:0] cache_0_s2_translator_avalon_universal_slave_0_agent_m0_address;                                          // cache_0_s2_translator_avalon_universal_slave_0_agent:m0_address -> cache_0_s2_translator:uav_address
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_m0_write;                                            // cache_0_s2_translator_avalon_universal_slave_0_agent:m0_write -> cache_0_s2_translator:uav_write
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_m0_lock;                                             // cache_0_s2_translator_avalon_universal_slave_0_agent:m0_lock -> cache_0_s2_translator:uav_lock
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_m0_read;                                             // cache_0_s2_translator_avalon_universal_slave_0_agent:m0_read -> cache_0_s2_translator:uav_read
	wire   [31:0] cache_0_s2_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // cache_0_s2_translator:uav_readdata -> cache_0_s2_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // cache_0_s2_translator:uav_readdatavalid -> cache_0_s2_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // cache_0_s2_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cache_0_s2_translator:uav_debugaccess
	wire    [3:0] cache_0_s2_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // cache_0_s2_translator_avalon_universal_slave_0_agent:m0_byteenable -> cache_0_s2_translator:uav_byteenable
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // cache_0_s2_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // cache_0_s2_translator_avalon_universal_slave_0_agent:rf_source_valid -> cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // cache_0_s2_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // cache_0_s2_translator_avalon_universal_slave_0_agent:rf_source_data -> cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cache_0_s2_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cache_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cache_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cache_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cache_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // cache_0_s2_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // cache_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // cache_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cache_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cache_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cache_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // cache_0_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_waitrequest;                          // distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_waitrequest -> distancecore_1_avalon_master_1_translator:uav_waitrequest
	wire    [2:0] distancecore_1_avalon_master_1_translator_avalon_universal_master_0_burstcount;                           // distancecore_1_avalon_master_1_translator:uav_burstcount -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] distancecore_1_avalon_master_1_translator_avalon_universal_master_0_writedata;                            // distancecore_1_avalon_master_1_translator:uav_writedata -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] distancecore_1_avalon_master_1_translator_avalon_universal_master_0_address;                              // distancecore_1_avalon_master_1_translator:uav_address -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_address
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_lock;                                 // distancecore_1_avalon_master_1_translator:uav_lock -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_lock
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_write;                                // distancecore_1_avalon_master_1_translator:uav_write -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_write
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_read;                                 // distancecore_1_avalon_master_1_translator:uav_read -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] distancecore_1_avalon_master_1_translator_avalon_universal_master_0_readdata;                             // distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_readdata -> distancecore_1_avalon_master_1_translator:uav_readdata
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_debugaccess;                          // distancecore_1_avalon_master_1_translator:uav_debugaccess -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] distancecore_1_avalon_master_1_translator_avalon_universal_master_0_byteenable;                           // distancecore_1_avalon_master_1_translator:uav_byteenable -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_byteenable
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_readdatavalid;                        // distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:av_readdatavalid -> distancecore_1_avalon_master_1_translator:uav_readdatavalid
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // cache_1_s2_translator:uav_waitrequest -> cache_1_s2_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cache_1_s2_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // cache_1_s2_translator_avalon_universal_slave_0_agent:m0_burstcount -> cache_1_s2_translator:uav_burstcount
	wire   [31:0] cache_1_s2_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // cache_1_s2_translator_avalon_universal_slave_0_agent:m0_writedata -> cache_1_s2_translator:uav_writedata
	wire   [15:0] cache_1_s2_translator_avalon_universal_slave_0_agent_m0_address;                                          // cache_1_s2_translator_avalon_universal_slave_0_agent:m0_address -> cache_1_s2_translator:uav_address
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_m0_write;                                            // cache_1_s2_translator_avalon_universal_slave_0_agent:m0_write -> cache_1_s2_translator:uav_write
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_m0_lock;                                             // cache_1_s2_translator_avalon_universal_slave_0_agent:m0_lock -> cache_1_s2_translator:uav_lock
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_m0_read;                                             // cache_1_s2_translator_avalon_universal_slave_0_agent:m0_read -> cache_1_s2_translator:uav_read
	wire   [31:0] cache_1_s2_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // cache_1_s2_translator:uav_readdata -> cache_1_s2_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // cache_1_s2_translator:uav_readdatavalid -> cache_1_s2_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // cache_1_s2_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cache_1_s2_translator:uav_debugaccess
	wire    [3:0] cache_1_s2_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // cache_1_s2_translator_avalon_universal_slave_0_agent:m0_byteenable -> cache_1_s2_translator:uav_byteenable
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // cache_1_s2_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // cache_1_s2_translator_avalon_universal_slave_0_agent:rf_source_valid -> cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // cache_1_s2_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // cache_1_s2_translator_avalon_universal_slave_0_agent:rf_source_data -> cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cache_1_s2_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cache_1_s2_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cache_1_s2_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cache_1_s2_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cache_1_s2_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // cache_1_s2_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // cache_1_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // cache_1_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cache_1_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cache_1_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cache_1_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // cache_1_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_waitrequest;                          // distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_waitrequest -> distancecore_2_avalon_master_1_translator:uav_waitrequest
	wire    [2:0] distancecore_2_avalon_master_1_translator_avalon_universal_master_0_burstcount;                           // distancecore_2_avalon_master_1_translator:uav_burstcount -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] distancecore_2_avalon_master_1_translator_avalon_universal_master_0_writedata;                            // distancecore_2_avalon_master_1_translator:uav_writedata -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_writedata
	wire   [15:0] distancecore_2_avalon_master_1_translator_avalon_universal_master_0_address;                              // distancecore_2_avalon_master_1_translator:uav_address -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_address
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_lock;                                 // distancecore_2_avalon_master_1_translator:uav_lock -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_lock
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_write;                                // distancecore_2_avalon_master_1_translator:uav_write -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_write
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_read;                                 // distancecore_2_avalon_master_1_translator:uav_read -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] distancecore_2_avalon_master_1_translator_avalon_universal_master_0_readdata;                             // distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_readdata -> distancecore_2_avalon_master_1_translator:uav_readdata
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_debugaccess;                          // distancecore_2_avalon_master_1_translator:uav_debugaccess -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] distancecore_2_avalon_master_1_translator_avalon_universal_master_0_byteenable;                           // distancecore_2_avalon_master_1_translator:uav_byteenable -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_byteenable
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_readdatavalid;                        // distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:av_readdatavalid -> distancecore_2_avalon_master_1_translator:uav_readdatavalid
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                      // cache_2_s2_translator:uav_waitrequest -> cache_2_s2_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cache_2_s2_translator_avalon_universal_slave_0_agent_m0_burstcount;                                       // cache_2_s2_translator_avalon_universal_slave_0_agent:m0_burstcount -> cache_2_s2_translator:uav_burstcount
	wire   [31:0] cache_2_s2_translator_avalon_universal_slave_0_agent_m0_writedata;                                        // cache_2_s2_translator_avalon_universal_slave_0_agent:m0_writedata -> cache_2_s2_translator:uav_writedata
	wire   [15:0] cache_2_s2_translator_avalon_universal_slave_0_agent_m0_address;                                          // cache_2_s2_translator_avalon_universal_slave_0_agent:m0_address -> cache_2_s2_translator:uav_address
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_m0_write;                                            // cache_2_s2_translator_avalon_universal_slave_0_agent:m0_write -> cache_2_s2_translator:uav_write
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_m0_lock;                                             // cache_2_s2_translator_avalon_universal_slave_0_agent:m0_lock -> cache_2_s2_translator:uav_lock
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_m0_read;                                             // cache_2_s2_translator_avalon_universal_slave_0_agent:m0_read -> cache_2_s2_translator:uav_read
	wire   [31:0] cache_2_s2_translator_avalon_universal_slave_0_agent_m0_readdata;                                         // cache_2_s2_translator:uav_readdata -> cache_2_s2_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                    // cache_2_s2_translator:uav_readdatavalid -> cache_2_s2_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                      // cache_2_s2_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cache_2_s2_translator:uav_debugaccess
	wire    [3:0] cache_2_s2_translator_avalon_universal_slave_0_agent_m0_byteenable;                                       // cache_2_s2_translator_avalon_universal_slave_0_agent:m0_byteenable -> cache_2_s2_translator:uav_byteenable
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                               // cache_2_s2_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_valid;                                     // cache_2_s2_translator_avalon_universal_slave_0_agent:rf_source_valid -> cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                             // cache_2_s2_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [85:0] cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_data;                                      // cache_2_s2_translator_avalon_universal_slave_0_agent:rf_source_data -> cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_ready;                                     // cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cache_2_s2_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                            // cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cache_2_s2_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                  // cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cache_2_s2_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                          // cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cache_2_s2_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [85:0] cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                   // cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cache_2_s2_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                  // cache_2_s2_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                // cache_2_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [31:0] cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                 // cache_2_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                // cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cache_2_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                // cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cache_2_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                 // cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cache_2_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                // cache_2_s2_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                             // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [102:0] cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                              // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router:sink_ready -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                    // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [102:0] cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                     // cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router_001:sink_ready -> cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                // dma_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_valid;                                      // dma_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                              // dma_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [102:0] dma_read_master_translator_avalon_universal_master_0_agent_cp_data;                                       // dma_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          dma_read_master_translator_avalon_universal_master_0_agent_cp_ready;                                      // addr_router_002:sink_ready -> dma_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [102:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [102:0] dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                                 // dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_001:sink_ready -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [102:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_002:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                              // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [102:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                               // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_003:sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                          // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire   [84:0] usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                           // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_004:sink_ready -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [102:0] sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_005:sink_ready -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [102:0] performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [102:0] ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                 // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_007:sink_ready -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                           // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [102:0] endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                            // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_008:sink_ready -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                              // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [102:0] fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                               // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_009:sink_ready -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                              // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [102:0] fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                               // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_010:sink_ready -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                               // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [102:0] ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_011:sink_ready -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                               // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [102:0] ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_012:sink_ready -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                             // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [102:0] emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                              // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_013:sink_ready -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                             // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [102:0] emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                              // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_014:sink_ready -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                           // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [102:0] endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                            // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_015:sink_ready -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                            // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [102:0] baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                             // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_016:sink_ready -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                          // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [102:0] skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                           // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_017:sink_ready -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                           // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [102:0] knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                            // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_018:sink_ready -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                             // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [102:0] emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                              // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_019:sink_ready -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                           // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [102:0] endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                            // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_020:sink_ready -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                              // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [102:0] fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                               // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire          fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_021:sink_ready -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                               // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	wire  [102:0] ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	wire          ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_022:sink_ready -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                               // dma_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_valid;                                     // dma_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                             // dma_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire   [86:0] dma_write_master_translator_avalon_universal_master_0_agent_cp_data;                                      // dma_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          dma_write_master_translator_avalon_universal_master_0_agent_cp_ready;                                     // addr_router_003:sink_ready -> dma_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                         // distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire   [86:0] distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                          // distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router_004:sink_ready -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                         // distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire   [86:0] distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                          // distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router_005:sink_ready -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                         // distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire   [86:0] distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                          // distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire          distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router_006:sink_ready -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // cache_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // cache_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // cache_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	wire   [86:0] cache_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // cache_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	wire          cache_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_023:sink_ready -> cache_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // cache_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // cache_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // cache_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	wire   [86:0] cache_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // cache_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	wire          cache_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_024:sink_ready -> cache_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // cache_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                            // cache_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // cache_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	wire   [86:0] cache_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                             // cache_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	wire          cache_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_025:sink_ready -> cache_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid;                       // distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket;               // distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire   [84:0] distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data;                        // distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire          distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_007:sink_ready -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:cp_ready
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // cache_0_s2_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rp_valid;                                            // cache_0_s2_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // cache_0_s2_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	wire   [84:0] cache_0_s2_translator_avalon_universal_slave_0_agent_rp_data;                                             // cache_0_s2_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	wire          cache_0_s2_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_026:sink_ready -> cache_0_s2_translator_avalon_universal_slave_0_agent:rp_ready
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid;                       // distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket;               // distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	wire   [84:0] distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data;                        // distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	wire          distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_008:sink_ready -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:cp_ready
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // cache_1_s2_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_027:sink_endofpacket
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rp_valid;                                            // cache_1_s2_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_027:sink_valid
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // cache_1_s2_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_027:sink_startofpacket
	wire   [84:0] cache_1_s2_translator_avalon_universal_slave_0_agent_rp_data;                                             // cache_1_s2_translator_avalon_universal_slave_0_agent:rp_data -> id_router_027:sink_data
	wire          cache_1_s2_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_027:sink_ready -> cache_1_s2_translator_avalon_universal_slave_0_agent:rp_ready
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_009:sink_endofpacket
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid;                       // distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_009:sink_valid
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket;               // distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_009:sink_startofpacket
	wire   [84:0] distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data;                        // distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:cp_data -> addr_router_009:sink_data
	wire          distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_009:sink_ready -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:cp_ready
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                      // cache_2_s2_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_028:sink_endofpacket
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rp_valid;                                            // cache_2_s2_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_028:sink_valid
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                    // cache_2_s2_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_028:sink_startofpacket
	wire   [84:0] cache_2_s2_translator_avalon_universal_slave_0_agent_rp_data;                                             // cache_2_s2_translator_avalon_universal_slave_0_agent:rp_data -> id_router_028:sink_data
	wire          cache_2_s2_translator_avalon_universal_slave_0_agent_rp_ready;                                            // id_router_028:sink_ready -> cache_2_s2_translator_avalon_universal_slave_0_agent:rp_ready
	wire          burst_adapter_source0_endofpacket;                                                                        // burst_adapter:source0_endofpacket -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                              // burst_adapter:source0_valid -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                      // burst_adapter:source0_startofpacket -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] burst_adapter_source0_data;                                                                               // burst_adapter:source0_data -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                              // usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [22:0] burst_adapter_source0_channel;                                                                            // burst_adapter:source0_channel -> usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                           // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, cache_0:reset, cache_0:reset2, cache_0_s1_translator:reset, cache_0_s1_translator_avalon_universal_slave_0_agent:reset, cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cache_0_s2_translator:reset, cache_0_s2_translator_avalon_universal_slave_0_agent:reset, cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cache_1:reset, cache_1:reset2, cache_1_s1_translator:reset, cache_1_s1_translator_avalon_universal_slave_0_agent:reset, cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cache_1_s2_translator:reset, cache_1_s2_translator_avalon_universal_slave_0_agent:reset, cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cache_2:reset, cache_2:reset2, cache_2_s1_translator:reset, cache_2_s1_translator_avalon_universal_slave_0_agent:reset, cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cache_2_s2_translator:reset, cache_2_s2_translator_avalon_universal_slave_0_agent:reset, cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_023:reset, cmd_xbar_mux_024:reset, cmd_xbar_mux_025:reset, cpu_0:reset_n, cpu_0_data_master_translator:reset, cpu_0_data_master_translator_avalon_universal_master_0_agent:reset, cpu_0_instruction_master_translator:reset, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:in_reset, crosser_007:in_reset, crosser_008:in_reset, crosser_009:in_reset, crosser_010:in_reset, crosser_011:in_reset, crosser_012:in_reset, crosser_013:in_reset, crosser_014:in_reset, crosser_015:in_reset, crosser_016:in_reset, crosser_017:out_reset, crosser_018:out_reset, crosser_019:out_reset, crosser_020:out_reset, crosser_021:out_reset, crosser_022:out_reset, crosser_023:out_reset, crosser_024:out_reset, crosser_025:out_reset, crosser_026:out_reset, crosser_027:out_reset, crosser_028:out_reset, crosser_029:out_reset, crosser_030:out_reset, crosser_031:out_reset, crosser_032:out_reset, crosser_033:out_reset, crosser_034:out_reset, crosser_035:out_reset, crosser_036:out_reset, crosser_037:in_reset, crosser_038:in_reset, crosser_039:in_reset, crosser_040:out_reset, crosser_041:in_reset, crosser_042:out_reset, crosser_043:in_reset, crosser_044:out_reset, crosser_045:in_reset, dma:system_reset_n, dma_control_port_slave_translator:reset, dma_control_port_slave_translator_avalon_universal_slave_0_agent:reset, dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_read_master_translator:reset, dma_read_master_translator_avalon_universal_master_0_agent:reset, dma_write_master_translator:reset, dma_write_master_translator_avalon_universal_master_0_agent:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_005:reset, id_router_006:reset, id_router_023:reset, id_router_024:reset, id_router_025:reset, id_router_026:reset, id_router_027:reset, id_router_028:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, performance_counter_0:reset_n, performance_counter_0_control_slave_translator:reset, performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_0:reset_n, pio_0_s1_translator:reset, pio_0_s1_translator_avalon_universal_slave_0_agent:reset, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rsp_xbar_demux_027:reset, rsp_xbar_demux_028:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_003:reset, sdram_controller:reset_n, sdram_controller_s1_translator:reset, sdram_controller_s1_translator_avalon_universal_slave_0_agent:reset, sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_001_reset_out_reset;                                                                       // rst_controller_001:reset_out -> [burst_adapter:reset, crosser:out_reset, crosser_017:in_reset, id_router_004:reset, rsp_xbar_demux_004:reset, usbFIFOCtrl_0:reset_n, usbFIFOCtrl_0_avalon_slave_0_translator:reset, usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, usbFIFOCtrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire          rst_controller_002_reset_out_reset;                                                                       // rst_controller_002:reset_out -> altpll_0:reset
	wire          rst_controller_003_reset_out_reset;                                                                       // rst_controller_003:reset_out -> [EndTSetReg_0:reset_n, EndTSetReg_0_avalon_slave_0_translator:reset, EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, EndTSetReg_1:reset_n, EndTSetReg_1_avalon_slave_0_translator:reset, EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, EndTSetReg_2:reset_n, EndTSetReg_2_avalon_slave_0_translator:reset, EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FullReg_0:reset_n, FullReg_0_avalon_slave_0_translator:reset, FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FullReg_1:reset_n, FullReg_1_avalon_slave_0_translator:reset, FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, FullReg_2:reset_n, FullReg_2_avalon_slave_0_translator:reset, FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, NDimReg:reset_n, NDimReg_avalon_slave_0_translator:reset, NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, NTrReg_0:reset_n, NTrReg_0_avalon_slave_0_translator:reset, NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, NTrReg_1:reset_n, NTrReg_1_avalon_slave_0_translator:reset, NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, NTrReg_2:reset_n, NTrReg_2_avalon_slave_0_translator:reset, NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router_004:reset, addr_router_005:reset, addr_router_006:reset, addr_router_007:reset, addr_router_008:reset, addr_router_009:reset, baseqaddr_0:reset_n, baseqaddr_0_avalon_slave_0_translator:reset, baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_007:reset, cmd_xbar_demux_008:reset, cmd_xbar_demux_009:reset, crosser_001:out_reset, crosser_002:out_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:out_reset, crosser_007:out_reset, crosser_008:out_reset, crosser_009:out_reset, crosser_010:out_reset, crosser_011:out_reset, crosser_012:out_reset, crosser_013:out_reset, crosser_014:out_reset, crosser_015:out_reset, crosser_016:out_reset, crosser_018:in_reset, crosser_019:in_reset, crosser_020:in_reset, crosser_021:in_reset, crosser_022:in_reset, crosser_023:in_reset, crosser_024:in_reset, crosser_025:in_reset, crosser_026:in_reset, crosser_027:in_reset, crosser_028:in_reset, crosser_029:in_reset, crosser_030:in_reset, crosser_031:in_reset, crosser_032:in_reset, crosser_033:in_reset, crosser_034:in_reset, crosser_035:in_reset, crosser_036:in_reset, crosser_037:out_reset, crosser_038:out_reset, crosser_039:out_reset, crosser_040:in_reset, crosser_041:out_reset, crosser_042:in_reset, crosser_043:out_reset, crosser_044:in_reset, crosser_045:out_reset, distancecore_0:reset_n, distancecore_0_avalon_master_1_translator:reset, distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:reset, distancecore_0_avalon_master_translator:reset, distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:reset, distancecore_1:reset_n, distancecore_1_avalon_master_1_translator:reset, distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:reset, distancecore_1_avalon_master_translator:reset, distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:reset, distancecore_2:reset_n, distancecore_2_avalon_master_1_translator:reset, distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:reset, distancecore_2_avalon_master_translator:reset, distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:reset, emptyreg_0:reset_n, emptyreg_0_avalon_slave_0_translator:reset, emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, emptyreg_1:reset_n, emptyreg_1_avalon_slave_0_translator:reset, emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, emptyreg_2:reset_n, emptyreg_2_avalon_slave_0_translator:reset, emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, knnclasscore:Reset, knnclasscore_avalon_slave_0_translator:reset, knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, skipaddrreg_0:reset_n, skipaddrreg_0_avalon_slave_0_translator:reset, skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_004_reset_out_reset;                                                                       // rst_controller_004:reset_out -> altpll_1:reset
	wire          cmd_xbar_demux_src0_endofpacket;                                                                          // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                        // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src0_data;                                                                                 // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [22:0] cmd_xbar_demux_src0_channel;                                                                              // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                          // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                        // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_src1_data;                                                                                 // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [22:0] cmd_xbar_demux_src1_channel;                                                                              // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                      // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                            // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                    // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src0_data;                                                                             // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [22:0] cmd_xbar_demux_001_src0_channel;                                                                          // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                            // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                      // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                            // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                    // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src1_data;                                                                             // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [22:0] cmd_xbar_demux_001_src1_channel;                                                                          // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                            // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                      // cmd_xbar_demux_001:src2_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                            // cmd_xbar_demux_001:src2_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                    // cmd_xbar_demux_001:src2_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src2_data;                                                                             // cmd_xbar_demux_001:src2_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src2_channel;                                                                          // cmd_xbar_demux_001:src2_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                      // cmd_xbar_demux_001:src3_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                            // cmd_xbar_demux_001:src3_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                    // cmd_xbar_demux_001:src3_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src3_data;                                                                             // cmd_xbar_demux_001:src3_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src3_channel;                                                                          // cmd_xbar_demux_001:src3_channel -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                      // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                            // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                    // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src5_data;                                                                             // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [22:0] cmd_xbar_demux_001_src5_channel;                                                                          // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                            // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux_001:src5_ready
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                      // cmd_xbar_demux_001:src6_endofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                            // cmd_xbar_demux_001:src6_valid -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                    // cmd_xbar_demux_001:src6_startofpacket -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src6_data;                                                                             // cmd_xbar_demux_001:src6_data -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_demux_001_src6_channel;                                                                          // cmd_xbar_demux_001:src6_channel -> performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                      // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                            // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                    // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [102:0] cmd_xbar_demux_002_src0_data;                                                                             // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_005:sink1_data
	wire   [22:0] cmd_xbar_demux_002_src0_channel;                                                                          // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                            // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                          // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                        // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [102:0] rsp_xbar_demux_src0_data;                                                                                 // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [22:0] rsp_xbar_demux_src0_channel;                                                                              // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                          // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                        // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [102:0] rsp_xbar_demux_src1_data;                                                                                 // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [22:0] rsp_xbar_demux_src1_channel;                                                                              // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                      // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                            // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                    // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [102:0] rsp_xbar_demux_001_src0_data;                                                                             // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [22:0] rsp_xbar_demux_001_src0_channel;                                                                          // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                            // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                      // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                            // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                    // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [102:0] rsp_xbar_demux_001_src1_data;                                                                             // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [22:0] rsp_xbar_demux_001_src1_channel;                                                                          // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                            // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                      // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                            // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                    // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [102:0] rsp_xbar_demux_002_src0_data;                                                                             // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [22:0] rsp_xbar_demux_002_src0_channel;                                                                          // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                            // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                      // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                            // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                    // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [102:0] rsp_xbar_demux_003_src0_data;                                                                             // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [22:0] rsp_xbar_demux_003_src0_channel;                                                                          // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                            // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                      // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                            // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                    // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [102:0] rsp_xbar_demux_005_src0_data;                                                                             // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [22:0] rsp_xbar_demux_005_src0_channel;                                                                          // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                            // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                      // rsp_xbar_demux_005:src1_endofpacket -> dma_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                            // rsp_xbar_demux_005:src1_valid -> dma_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                    // rsp_xbar_demux_005:src1_startofpacket -> dma_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_demux_005_src1_data;                                                                             // rsp_xbar_demux_005:src1_data -> dma_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [22:0] rsp_xbar_demux_005_src1_channel;                                                                          // rsp_xbar_demux_005:src1_channel -> dma_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                      // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                            // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                    // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [102:0] rsp_xbar_demux_006_src0_data;                                                                             // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [22:0] rsp_xbar_demux_006_src0_channel;                                                                          // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                            // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          addr_router_src_endofpacket;                                                                              // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                                    // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                            // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [102:0] addr_router_src_data;                                                                                     // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [22:0] addr_router_src_channel;                                                                                  // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                                    // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                             // rsp_xbar_mux:src_endofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                   // rsp_xbar_mux:src_valid -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                           // rsp_xbar_mux:src_startofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_mux_src_data;                                                                                    // rsp_xbar_mux:src_data -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [22:0] rsp_xbar_mux_src_channel;                                                                                 // rsp_xbar_mux:src_channel -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                                   // cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                          // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                        // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [102:0] addr_router_001_src_data;                                                                                 // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [22:0] addr_router_001_src_channel;                                                                              // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                                // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                         // rsp_xbar_mux_001:src_endofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                               // rsp_xbar_mux_001:src_valid -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                       // rsp_xbar_mux_001:src_startofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [102:0] rsp_xbar_mux_001_src_data;                                                                                // rsp_xbar_mux_001:src_data -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [22:0] rsp_xbar_mux_001_src_channel;                                                                             // rsp_xbar_mux_001:src_channel -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                               // cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                          // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                        // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [102:0] addr_router_002_src_data;                                                                                 // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [22:0] addr_router_002_src_channel;                                                                              // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_005_src1_ready;                                                                            // dma_read_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_005:src1_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                             // cmd_xbar_mux:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                   // cmd_xbar_mux:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                           // cmd_xbar_mux:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_src_data;                                                                                    // cmd_xbar_mux:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_mux_src_channel;                                                                                 // cmd_xbar_mux:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                      // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                              // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [102:0] id_router_src_data;                                                                                       // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [22:0] id_router_src_channel;                                                                                    // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                      // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                         // cmd_xbar_mux_001:src_endofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                               // cmd_xbar_mux_001:src_valid -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                       // cmd_xbar_mux_001:src_startofpacket -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_001_src_data;                                                                                // cmd_xbar_mux_001:src_data -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_mux_001_src_channel;                                                                             // cmd_xbar_mux_001:src_channel -> dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                               // dma_control_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                            // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                  // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                          // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [102:0] id_router_001_src_data;                                                                                   // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [22:0] id_router_001_src_channel;                                                                                // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                  // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_001_src2_ready;                                                                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire          id_router_002_src_endofpacket;                                                                            // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                  // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                          // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [102:0] id_router_002_src_data;                                                                                   // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [22:0] id_router_002_src_channel;                                                                                // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                  // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_demux_001_src3_ready;                                                                            // pio_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire          id_router_003_src_endofpacket;                                                                            // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                  // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                          // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [102:0] id_router_003_src_data;                                                                                   // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [22:0] id_router_003_src_channel;                                                                                // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                  // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                         // cmd_xbar_mux_005:src_endofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                               // cmd_xbar_mux_005:src_valid -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                       // cmd_xbar_mux_005:src_startofpacket -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] cmd_xbar_mux_005_src_data;                                                                                // cmd_xbar_mux_005:src_data -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] cmd_xbar_mux_005_src_channel;                                                                             // cmd_xbar_mux_005:src_channel -> sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                               // sdram_controller_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                            // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                  // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                          // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [102:0] id_router_005_src_data;                                                                                   // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [22:0] id_router_005_src_channel;                                                                                // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                  // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                            // performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                            // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                  // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                          // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [102:0] id_router_006_src_data;                                                                                   // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [22:0] id_router_006_src_channel;                                                                                // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                  // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          crosser_001_out_ready;                                                                                    // NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	wire          id_router_007_src_endofpacket;                                                                            // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                  // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                          // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [102:0] id_router_007_src_data;                                                                                   // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [22:0] id_router_007_src_channel;                                                                                // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                  // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          crosser_002_out_ready;                                                                                    // EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_002:out_ready
	wire          id_router_008_src_endofpacket;                                                                            // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                  // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                          // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [102:0] id_router_008_src_data;                                                                                   // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [22:0] id_router_008_src_channel;                                                                                // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                  // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          crosser_003_out_ready;                                                                                    // FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_003:out_ready
	wire          id_router_009_src_endofpacket;                                                                            // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                  // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                          // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [102:0] id_router_009_src_data;                                                                                   // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [22:0] id_router_009_src_channel;                                                                                // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                  // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          crosser_004_out_ready;                                                                                    // FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_004:out_ready
	wire          id_router_010_src_endofpacket;                                                                            // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                  // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                          // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [102:0] id_router_010_src_data;                                                                                   // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [22:0] id_router_010_src_channel;                                                                                // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                  // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          crosser_005_out_ready;                                                                                    // NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_005:out_ready
	wire          id_router_011_src_endofpacket;                                                                            // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                  // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                          // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [102:0] id_router_011_src_data;                                                                                   // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [22:0] id_router_011_src_channel;                                                                                // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                  // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          crosser_006_out_ready;                                                                                    // NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_006:out_ready
	wire          id_router_012_src_endofpacket;                                                                            // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                  // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                          // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [102:0] id_router_012_src_data;                                                                                   // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [22:0] id_router_012_src_channel;                                                                                // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                  // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          crosser_007_out_ready;                                                                                    // emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_007:out_ready
	wire          id_router_013_src_endofpacket;                                                                            // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                  // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                          // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [102:0] id_router_013_src_data;                                                                                   // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [22:0] id_router_013_src_channel;                                                                                // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                  // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          crosser_008_out_ready;                                                                                    // emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_008:out_ready
	wire          id_router_014_src_endofpacket;                                                                            // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                  // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                          // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [102:0] id_router_014_src_data;                                                                                   // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [22:0] id_router_014_src_channel;                                                                                // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                  // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          crosser_009_out_ready;                                                                                    // EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_009:out_ready
	wire          id_router_015_src_endofpacket;                                                                            // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                  // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                          // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [102:0] id_router_015_src_data;                                                                                   // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [22:0] id_router_015_src_channel;                                                                                // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                  // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          crosser_010_out_ready;                                                                                    // baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_010:out_ready
	wire          id_router_016_src_endofpacket;                                                                            // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                  // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                          // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [102:0] id_router_016_src_data;                                                                                   // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [22:0] id_router_016_src_channel;                                                                                // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                  // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          crosser_011_out_ready;                                                                                    // skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_011:out_ready
	wire          id_router_017_src_endofpacket;                                                                            // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                  // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                          // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [102:0] id_router_017_src_data;                                                                                   // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [22:0] id_router_017_src_channel;                                                                                // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                  // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          crosser_012_out_ready;                                                                                    // knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_012:out_ready
	wire          id_router_018_src_endofpacket;                                                                            // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                  // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                          // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [102:0] id_router_018_src_data;                                                                                   // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [22:0] id_router_018_src_channel;                                                                                // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                  // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          crosser_013_out_ready;                                                                                    // emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_013:out_ready
	wire          id_router_019_src_endofpacket;                                                                            // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          id_router_019_src_valid;                                                                                  // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire          id_router_019_src_startofpacket;                                                                          // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [102:0] id_router_019_src_data;                                                                                   // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire   [22:0] id_router_019_src_channel;                                                                                // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire          id_router_019_src_ready;                                                                                  // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire          crosser_014_out_ready;                                                                                    // EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_014:out_ready
	wire          id_router_020_src_endofpacket;                                                                            // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          id_router_020_src_valid;                                                                                  // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire          id_router_020_src_startofpacket;                                                                          // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [102:0] id_router_020_src_data;                                                                                   // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire   [22:0] id_router_020_src_channel;                                                                                // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire          id_router_020_src_ready;                                                                                  // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire          crosser_015_out_ready;                                                                                    // FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_015:out_ready
	wire          id_router_021_src_endofpacket;                                                                            // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire          id_router_021_src_valid;                                                                                  // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire          id_router_021_src_startofpacket;                                                                          // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [102:0] id_router_021_src_data;                                                                                   // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire   [22:0] id_router_021_src_channel;                                                                                // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire          id_router_021_src_ready;                                                                                  // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire          crosser_016_out_ready;                                                                                    // NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_016:out_ready
	wire          id_router_022_src_endofpacket;                                                                            // id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	wire          id_router_022_src_valid;                                                                                  // id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	wire          id_router_022_src_startofpacket;                                                                          // id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	wire  [102:0] id_router_022_src_data;                                                                                   // id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	wire   [22:0] id_router_022_src_channel;                                                                                // id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	wire          id_router_022_src_ready;                                                                                  // rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                      // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_023:sink0_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                            // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_023:sink0_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                    // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_023:sink0_startofpacket
	wire   [86:0] cmd_xbar_demux_003_src0_data;                                                                             // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_023:sink0_data
	wire    [3:0] cmd_xbar_demux_003_src0_channel;                                                                          // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_023:sink0_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                            // cmd_xbar_mux_023:sink0_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                                      // cmd_xbar_demux_003:src1_endofpacket -> cmd_xbar_mux_024:sink0_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                            // cmd_xbar_demux_003:src1_valid -> cmd_xbar_mux_024:sink0_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                                    // cmd_xbar_demux_003:src1_startofpacket -> cmd_xbar_mux_024:sink0_startofpacket
	wire   [86:0] cmd_xbar_demux_003_src1_data;                                                                             // cmd_xbar_demux_003:src1_data -> cmd_xbar_mux_024:sink0_data
	wire    [3:0] cmd_xbar_demux_003_src1_channel;                                                                          // cmd_xbar_demux_003:src1_channel -> cmd_xbar_mux_024:sink0_channel
	wire          cmd_xbar_demux_003_src1_ready;                                                                            // cmd_xbar_mux_024:sink0_ready -> cmd_xbar_demux_003:src1_ready
	wire          cmd_xbar_demux_003_src2_endofpacket;                                                                      // cmd_xbar_demux_003:src2_endofpacket -> cmd_xbar_mux_025:sink0_endofpacket
	wire          cmd_xbar_demux_003_src2_valid;                                                                            // cmd_xbar_demux_003:src2_valid -> cmd_xbar_mux_025:sink0_valid
	wire          cmd_xbar_demux_003_src2_startofpacket;                                                                    // cmd_xbar_demux_003:src2_startofpacket -> cmd_xbar_mux_025:sink0_startofpacket
	wire   [86:0] cmd_xbar_demux_003_src2_data;                                                                             // cmd_xbar_demux_003:src2_data -> cmd_xbar_mux_025:sink0_data
	wire    [3:0] cmd_xbar_demux_003_src2_channel;                                                                          // cmd_xbar_demux_003:src2_channel -> cmd_xbar_mux_025:sink0_channel
	wire          cmd_xbar_demux_003_src2_ready;                                                                            // cmd_xbar_mux_025:sink0_ready -> cmd_xbar_demux_003:src2_ready
	wire          rsp_xbar_demux_023_src0_endofpacket;                                                                      // rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_023_src0_valid;                                                                            // rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_023_src0_startofpacket;                                                                    // rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire   [86:0] rsp_xbar_demux_023_src0_data;                                                                             // rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_003:sink0_data
	wire    [3:0] rsp_xbar_demux_023_src0_channel;                                                                          // rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_023_src0_ready;                                                                            // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_023:src0_ready
	wire          rsp_xbar_demux_024_src0_endofpacket;                                                                      // rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_024_src0_valid;                                                                            // rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_024_src0_startofpacket;                                                                    // rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire   [86:0] rsp_xbar_demux_024_src0_data;                                                                             // rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_003:sink1_data
	wire    [3:0] rsp_xbar_demux_024_src0_channel;                                                                          // rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_024_src0_ready;                                                                            // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_024:src0_ready
	wire          rsp_xbar_demux_025_src0_endofpacket;                                                                      // rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_003:sink2_endofpacket
	wire          rsp_xbar_demux_025_src0_valid;                                                                            // rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_003:sink2_valid
	wire          rsp_xbar_demux_025_src0_startofpacket;                                                                    // rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_003:sink2_startofpacket
	wire   [86:0] rsp_xbar_demux_025_src0_data;                                                                             // rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_003:sink2_data
	wire    [3:0] rsp_xbar_demux_025_src0_channel;                                                                          // rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_003:sink2_channel
	wire          rsp_xbar_demux_025_src0_ready;                                                                            // rsp_xbar_mux_003:sink2_ready -> rsp_xbar_demux_025:src0_ready
	wire          addr_router_003_src_endofpacket;                                                                          // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                                // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                        // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire   [86:0] addr_router_003_src_data;                                                                                 // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire    [3:0] addr_router_003_src_channel;                                                                              // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                                // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                         // rsp_xbar_mux_003:src_endofpacket -> dma_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                               // rsp_xbar_mux_003:src_valid -> dma_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                                       // rsp_xbar_mux_003:src_startofpacket -> dma_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [86:0] rsp_xbar_mux_003_src_data;                                                                                // rsp_xbar_mux_003:src_data -> dma_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] rsp_xbar_mux_003_src_channel;                                                                             // rsp_xbar_mux_003:src_channel -> dma_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                               // dma_write_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_003:src_ready
	wire          addr_router_004_src_endofpacket;                                                                          // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                                // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                        // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire   [86:0] addr_router_004_src_data;                                                                                 // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire    [3:0] addr_router_004_src_channel;                                                                              // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                                // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          crosser_039_out_ready;                                                                                    // distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> crosser_039:out_ready
	wire          addr_router_005_src_endofpacket;                                                                          // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          addr_router_005_src_valid;                                                                                // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire          addr_router_005_src_startofpacket;                                                                        // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire   [86:0] addr_router_005_src_data;                                                                                 // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire    [3:0] addr_router_005_src_channel;                                                                              // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire          addr_router_005_src_ready;                                                                                // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire          crosser_038_out_ready;                                                                                    // distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> crosser_038:out_ready
	wire          addr_router_006_src_endofpacket;                                                                          // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire          addr_router_006_src_valid;                                                                                // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire          addr_router_006_src_startofpacket;                                                                        // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire   [86:0] addr_router_006_src_data;                                                                                 // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire    [3:0] addr_router_006_src_channel;                                                                              // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire          addr_router_006_src_ready;                                                                                // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire          crosser_037_out_ready;                                                                                    // distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> crosser_037:out_ready
	wire          cmd_xbar_mux_023_src_endofpacket;                                                                         // cmd_xbar_mux_023:src_endofpacket -> cache_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_023_src_valid;                                                                               // cmd_xbar_mux_023:src_valid -> cache_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_023_src_startofpacket;                                                                       // cmd_xbar_mux_023:src_startofpacket -> cache_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [86:0] cmd_xbar_mux_023_src_data;                                                                                // cmd_xbar_mux_023:src_data -> cache_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_mux_023_src_channel;                                                                             // cmd_xbar_mux_023:src_channel -> cache_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_023_src_ready;                                                                               // cache_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_023:src_ready
	wire          id_router_023_src_endofpacket;                                                                            // id_router_023:src_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	wire          id_router_023_src_valid;                                                                                  // id_router_023:src_valid -> rsp_xbar_demux_023:sink_valid
	wire          id_router_023_src_startofpacket;                                                                          // id_router_023:src_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	wire   [86:0] id_router_023_src_data;                                                                                   // id_router_023:src_data -> rsp_xbar_demux_023:sink_data
	wire    [3:0] id_router_023_src_channel;                                                                                // id_router_023:src_channel -> rsp_xbar_demux_023:sink_channel
	wire          id_router_023_src_ready;                                                                                  // rsp_xbar_demux_023:sink_ready -> id_router_023:src_ready
	wire          cmd_xbar_mux_024_src_endofpacket;                                                                         // cmd_xbar_mux_024:src_endofpacket -> cache_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_024_src_valid;                                                                               // cmd_xbar_mux_024:src_valid -> cache_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_024_src_startofpacket;                                                                       // cmd_xbar_mux_024:src_startofpacket -> cache_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [86:0] cmd_xbar_mux_024_src_data;                                                                                // cmd_xbar_mux_024:src_data -> cache_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_mux_024_src_channel;                                                                             // cmd_xbar_mux_024:src_channel -> cache_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_024_src_ready;                                                                               // cache_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_024:src_ready
	wire          id_router_024_src_endofpacket;                                                                            // id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	wire          id_router_024_src_valid;                                                                                  // id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	wire          id_router_024_src_startofpacket;                                                                          // id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	wire   [86:0] id_router_024_src_data;                                                                                   // id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	wire    [3:0] id_router_024_src_channel;                                                                                // id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	wire          id_router_024_src_ready;                                                                                  // rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	wire          cmd_xbar_mux_025_src_endofpacket;                                                                         // cmd_xbar_mux_025:src_endofpacket -> cache_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_025_src_valid;                                                                               // cmd_xbar_mux_025:src_valid -> cache_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_025_src_startofpacket;                                                                       // cmd_xbar_mux_025:src_startofpacket -> cache_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [86:0] cmd_xbar_mux_025_src_data;                                                                                // cmd_xbar_mux_025:src_data -> cache_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_mux_025_src_channel;                                                                             // cmd_xbar_mux_025:src_channel -> cache_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_025_src_ready;                                                                               // cache_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_025:src_ready
	wire          id_router_025_src_endofpacket;                                                                            // id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	wire          id_router_025_src_valid;                                                                                  // id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	wire          id_router_025_src_startofpacket;                                                                          // id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	wire   [86:0] id_router_025_src_data;                                                                                   // id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	wire    [3:0] id_router_025_src_channel;                                                                                // id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	wire          id_router_025_src_ready;                                                                                  // rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	wire          addr_router_007_src_endofpacket;                                                                          // addr_router_007:src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire          addr_router_007_src_valid;                                                                                // addr_router_007:src_valid -> cmd_xbar_demux_007:sink_valid
	wire          addr_router_007_src_startofpacket;                                                                        // addr_router_007:src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire   [84:0] addr_router_007_src_data;                                                                                 // addr_router_007:src_data -> cmd_xbar_demux_007:sink_data
	wire    [0:0] addr_router_007_src_channel;                                                                              // addr_router_007:src_channel -> cmd_xbar_demux_007:sink_channel
	wire          addr_router_007_src_ready;                                                                                // cmd_xbar_demux_007:sink_ready -> addr_router_007:src_ready
	wire          crosser_041_out_ready;                                                                                    // distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:rp_ready -> crosser_041:out_ready
	wire          crosser_040_out_ready;                                                                                    // cache_0_s2_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_040:out_ready
	wire          id_router_026_src_endofpacket;                                                                            // id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	wire          id_router_026_src_valid;                                                                                  // id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	wire          id_router_026_src_startofpacket;                                                                          // id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	wire   [84:0] id_router_026_src_data;                                                                                   // id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	wire    [0:0] id_router_026_src_channel;                                                                                // id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	wire          id_router_026_src_ready;                                                                                  // rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	wire          addr_router_008_src_endofpacket;                                                                          // addr_router_008:src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	wire          addr_router_008_src_valid;                                                                                // addr_router_008:src_valid -> cmd_xbar_demux_008:sink_valid
	wire          addr_router_008_src_startofpacket;                                                                        // addr_router_008:src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	wire   [84:0] addr_router_008_src_data;                                                                                 // addr_router_008:src_data -> cmd_xbar_demux_008:sink_data
	wire    [0:0] addr_router_008_src_channel;                                                                              // addr_router_008:src_channel -> cmd_xbar_demux_008:sink_channel
	wire          addr_router_008_src_ready;                                                                                // cmd_xbar_demux_008:sink_ready -> addr_router_008:src_ready
	wire          crosser_043_out_ready;                                                                                    // distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:rp_ready -> crosser_043:out_ready
	wire          crosser_042_out_ready;                                                                                    // cache_1_s2_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_042:out_ready
	wire          id_router_027_src_endofpacket;                                                                            // id_router_027:src_endofpacket -> rsp_xbar_demux_027:sink_endofpacket
	wire          id_router_027_src_valid;                                                                                  // id_router_027:src_valid -> rsp_xbar_demux_027:sink_valid
	wire          id_router_027_src_startofpacket;                                                                          // id_router_027:src_startofpacket -> rsp_xbar_demux_027:sink_startofpacket
	wire   [84:0] id_router_027_src_data;                                                                                   // id_router_027:src_data -> rsp_xbar_demux_027:sink_data
	wire    [0:0] id_router_027_src_channel;                                                                                // id_router_027:src_channel -> rsp_xbar_demux_027:sink_channel
	wire          id_router_027_src_ready;                                                                                  // rsp_xbar_demux_027:sink_ready -> id_router_027:src_ready
	wire          addr_router_009_src_endofpacket;                                                                          // addr_router_009:src_endofpacket -> cmd_xbar_demux_009:sink_endofpacket
	wire          addr_router_009_src_valid;                                                                                // addr_router_009:src_valid -> cmd_xbar_demux_009:sink_valid
	wire          addr_router_009_src_startofpacket;                                                                        // addr_router_009:src_startofpacket -> cmd_xbar_demux_009:sink_startofpacket
	wire   [84:0] addr_router_009_src_data;                                                                                 // addr_router_009:src_data -> cmd_xbar_demux_009:sink_data
	wire    [0:0] addr_router_009_src_channel;                                                                              // addr_router_009:src_channel -> cmd_xbar_demux_009:sink_channel
	wire          addr_router_009_src_ready;                                                                                // cmd_xbar_demux_009:sink_ready -> addr_router_009:src_ready
	wire          crosser_045_out_ready;                                                                                    // distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:rp_ready -> crosser_045:out_ready
	wire          crosser_044_out_ready;                                                                                    // cache_2_s2_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_044:out_ready
	wire          id_router_028_src_endofpacket;                                                                            // id_router_028:src_endofpacket -> rsp_xbar_demux_028:sink_endofpacket
	wire          id_router_028_src_valid;                                                                                  // id_router_028:src_valid -> rsp_xbar_demux_028:sink_valid
	wire          id_router_028_src_startofpacket;                                                                          // id_router_028:src_startofpacket -> rsp_xbar_demux_028:sink_startofpacket
	wire   [84:0] id_router_028_src_data;                                                                                   // id_router_028:src_data -> rsp_xbar_demux_028:sink_data
	wire    [0:0] id_router_028_src_channel;                                                                                // id_router_028:src_channel -> rsp_xbar_demux_028:sink_channel
	wire          id_router_028_src_ready;                                                                                  // rsp_xbar_demux_028:sink_ready -> id_router_028:src_ready
	wire          crosser_out_ready;                                                                                        // width_adapter:in_ready -> crosser:out_ready
	wire          width_adapter_src_endofpacket;                                                                            // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                  // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                          // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [84:0] width_adapter_src_data;                                                                                   // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                                  // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [22:0] width_adapter_src_channel;                                                                                // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_004_src_endofpacket;                                                                            // id_router_004:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_004_src_valid;                                                                                  // id_router_004:src_valid -> width_adapter_001:in_valid
	wire          id_router_004_src_startofpacket;                                                                          // id_router_004:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [84:0] id_router_004_src_data;                                                                                   // id_router_004:src_data -> width_adapter_001:in_data
	wire   [22:0] id_router_004_src_channel;                                                                                // id_router_004:src_channel -> width_adapter_001:in_channel
	wire          id_router_004_src_ready;                                                                                  // width_adapter_001:in_ready -> id_router_004:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                        // width_adapter_001:out_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                              // width_adapter_001:out_valid -> rsp_xbar_demux_004:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                      // width_adapter_001:out_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [102:0] width_adapter_001_src_data;                                                                               // width_adapter_001:out_data -> rsp_xbar_demux_004:sink_data
	wire          width_adapter_001_src_ready;                                                                              // rsp_xbar_demux_004:sink_ready -> width_adapter_001:out_ready
	wire   [22:0] width_adapter_001_src_channel;                                                                            // width_adapter_001:out_channel -> rsp_xbar_demux_004:sink_channel
	wire          crosser_out_endofpacket;                                                                                  // crosser:out_endofpacket -> width_adapter:in_endofpacket
	wire          crosser_out_valid;                                                                                        // crosser:out_valid -> width_adapter:in_valid
	wire          crosser_out_startofpacket;                                                                                // crosser:out_startofpacket -> width_adapter:in_startofpacket
	wire  [102:0] crosser_out_data;                                                                                         // crosser:out_data -> width_adapter:in_data
	wire   [22:0] crosser_out_channel;                                                                                      // crosser:out_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                      // cmd_xbar_demux_001:src4_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                            // cmd_xbar_demux_001:src4_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                    // cmd_xbar_demux_001:src4_startofpacket -> crosser:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src4_data;                                                                             // cmd_xbar_demux_001:src4_data -> crosser:in_data
	wire   [22:0] cmd_xbar_demux_001_src4_channel;                                                                          // cmd_xbar_demux_001:src4_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                            // crosser:in_ready -> cmd_xbar_demux_001:src4_ready
	wire          crosser_001_out_endofpacket;                                                                              // crosser_001:out_endofpacket -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_001_out_valid;                                                                                    // crosser_001:out_valid -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_001_out_startofpacket;                                                                            // crosser_001:out_startofpacket -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_001_out_data;                                                                                     // crosser_001:out_data -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_001_out_channel;                                                                                  // crosser_001:out_channel -> NDimReg_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                      // cmd_xbar_demux_001:src7_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                            // cmd_xbar_demux_001:src7_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                    // cmd_xbar_demux_001:src7_startofpacket -> crosser_001:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src7_data;                                                                             // cmd_xbar_demux_001:src7_data -> crosser_001:in_data
	wire   [22:0] cmd_xbar_demux_001_src7_channel;                                                                          // cmd_xbar_demux_001:src7_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_001_src7_ready;                                                                            // crosser_001:in_ready -> cmd_xbar_demux_001:src7_ready
	wire          crosser_002_out_endofpacket;                                                                              // crosser_002:out_endofpacket -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_002_out_valid;                                                                                    // crosser_002:out_valid -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_002_out_startofpacket;                                                                            // crosser_002:out_startofpacket -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_002_out_data;                                                                                     // crosser_002:out_data -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_002_out_channel;                                                                                  // crosser_002:out_channel -> EndTSetReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                      // cmd_xbar_demux_001:src8_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                            // cmd_xbar_demux_001:src8_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                    // cmd_xbar_demux_001:src8_startofpacket -> crosser_002:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src8_data;                                                                             // cmd_xbar_demux_001:src8_data -> crosser_002:in_data
	wire   [22:0] cmd_xbar_demux_001_src8_channel;                                                                          // cmd_xbar_demux_001:src8_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_001_src8_ready;                                                                            // crosser_002:in_ready -> cmd_xbar_demux_001:src8_ready
	wire          crosser_003_out_endofpacket;                                                                              // crosser_003:out_endofpacket -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_003_out_valid;                                                                                    // crosser_003:out_valid -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_003_out_startofpacket;                                                                            // crosser_003:out_startofpacket -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_003_out_data;                                                                                     // crosser_003:out_data -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_003_out_channel;                                                                                  // crosser_003:out_channel -> FullReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                      // cmd_xbar_demux_001:src9_endofpacket -> crosser_003:in_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                            // cmd_xbar_demux_001:src9_valid -> crosser_003:in_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                    // cmd_xbar_demux_001:src9_startofpacket -> crosser_003:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src9_data;                                                                             // cmd_xbar_demux_001:src9_data -> crosser_003:in_data
	wire   [22:0] cmd_xbar_demux_001_src9_channel;                                                                          // cmd_xbar_demux_001:src9_channel -> crosser_003:in_channel
	wire          cmd_xbar_demux_001_src9_ready;                                                                            // crosser_003:in_ready -> cmd_xbar_demux_001:src9_ready
	wire          crosser_004_out_endofpacket;                                                                              // crosser_004:out_endofpacket -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_004_out_valid;                                                                                    // crosser_004:out_valid -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_004_out_startofpacket;                                                                            // crosser_004:out_startofpacket -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_004_out_data;                                                                                     // crosser_004:out_data -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_004_out_channel;                                                                                  // crosser_004:out_channel -> FullReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                     // cmd_xbar_demux_001:src10_endofpacket -> crosser_004:in_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                           // cmd_xbar_demux_001:src10_valid -> crosser_004:in_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                   // cmd_xbar_demux_001:src10_startofpacket -> crosser_004:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src10_data;                                                                            // cmd_xbar_demux_001:src10_data -> crosser_004:in_data
	wire   [22:0] cmd_xbar_demux_001_src10_channel;                                                                         // cmd_xbar_demux_001:src10_channel -> crosser_004:in_channel
	wire          cmd_xbar_demux_001_src10_ready;                                                                           // crosser_004:in_ready -> cmd_xbar_demux_001:src10_ready
	wire          crosser_005_out_endofpacket;                                                                              // crosser_005:out_endofpacket -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_005_out_valid;                                                                                    // crosser_005:out_valid -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_005_out_startofpacket;                                                                            // crosser_005:out_startofpacket -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_005_out_data;                                                                                     // crosser_005:out_data -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_005_out_channel;                                                                                  // crosser_005:out_channel -> NTrReg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                     // cmd_xbar_demux_001:src11_endofpacket -> crosser_005:in_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                           // cmd_xbar_demux_001:src11_valid -> crosser_005:in_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                   // cmd_xbar_demux_001:src11_startofpacket -> crosser_005:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src11_data;                                                                            // cmd_xbar_demux_001:src11_data -> crosser_005:in_data
	wire   [22:0] cmd_xbar_demux_001_src11_channel;                                                                         // cmd_xbar_demux_001:src11_channel -> crosser_005:in_channel
	wire          cmd_xbar_demux_001_src11_ready;                                                                           // crosser_005:in_ready -> cmd_xbar_demux_001:src11_ready
	wire          crosser_006_out_endofpacket;                                                                              // crosser_006:out_endofpacket -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_006_out_valid;                                                                                    // crosser_006:out_valid -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_006_out_startofpacket;                                                                            // crosser_006:out_startofpacket -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_006_out_data;                                                                                     // crosser_006:out_data -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_006_out_channel;                                                                                  // crosser_006:out_channel -> NTrReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                     // cmd_xbar_demux_001:src12_endofpacket -> crosser_006:in_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                           // cmd_xbar_demux_001:src12_valid -> crosser_006:in_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                   // cmd_xbar_demux_001:src12_startofpacket -> crosser_006:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src12_data;                                                                            // cmd_xbar_demux_001:src12_data -> crosser_006:in_data
	wire   [22:0] cmd_xbar_demux_001_src12_channel;                                                                         // cmd_xbar_demux_001:src12_channel -> crosser_006:in_channel
	wire          cmd_xbar_demux_001_src12_ready;                                                                           // crosser_006:in_ready -> cmd_xbar_demux_001:src12_ready
	wire          crosser_007_out_endofpacket;                                                                              // crosser_007:out_endofpacket -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_007_out_valid;                                                                                    // crosser_007:out_valid -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_007_out_startofpacket;                                                                            // crosser_007:out_startofpacket -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_007_out_data;                                                                                     // crosser_007:out_data -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_007_out_channel;                                                                                  // crosser_007:out_channel -> emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                     // cmd_xbar_demux_001:src13_endofpacket -> crosser_007:in_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                           // cmd_xbar_demux_001:src13_valid -> crosser_007:in_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                   // cmd_xbar_demux_001:src13_startofpacket -> crosser_007:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src13_data;                                                                            // cmd_xbar_demux_001:src13_data -> crosser_007:in_data
	wire   [22:0] cmd_xbar_demux_001_src13_channel;                                                                         // cmd_xbar_demux_001:src13_channel -> crosser_007:in_channel
	wire          cmd_xbar_demux_001_src13_ready;                                                                           // crosser_007:in_ready -> cmd_xbar_demux_001:src13_ready
	wire          crosser_008_out_endofpacket;                                                                              // crosser_008:out_endofpacket -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_008_out_valid;                                                                                    // crosser_008:out_valid -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_008_out_startofpacket;                                                                            // crosser_008:out_startofpacket -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_008_out_data;                                                                                     // crosser_008:out_data -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_008_out_channel;                                                                                  // crosser_008:out_channel -> emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                     // cmd_xbar_demux_001:src14_endofpacket -> crosser_008:in_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                           // cmd_xbar_demux_001:src14_valid -> crosser_008:in_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                   // cmd_xbar_demux_001:src14_startofpacket -> crosser_008:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src14_data;                                                                            // cmd_xbar_demux_001:src14_data -> crosser_008:in_data
	wire   [22:0] cmd_xbar_demux_001_src14_channel;                                                                         // cmd_xbar_demux_001:src14_channel -> crosser_008:in_channel
	wire          cmd_xbar_demux_001_src14_ready;                                                                           // crosser_008:in_ready -> cmd_xbar_demux_001:src14_ready
	wire          crosser_009_out_endofpacket;                                                                              // crosser_009:out_endofpacket -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_009_out_valid;                                                                                    // crosser_009:out_valid -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_009_out_startofpacket;                                                                            // crosser_009:out_startofpacket -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_009_out_data;                                                                                     // crosser_009:out_data -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_009_out_channel;                                                                                  // crosser_009:out_channel -> EndTSetReg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                     // cmd_xbar_demux_001:src15_endofpacket -> crosser_009:in_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                           // cmd_xbar_demux_001:src15_valid -> crosser_009:in_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                   // cmd_xbar_demux_001:src15_startofpacket -> crosser_009:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src15_data;                                                                            // cmd_xbar_demux_001:src15_data -> crosser_009:in_data
	wire   [22:0] cmd_xbar_demux_001_src15_channel;                                                                         // cmd_xbar_demux_001:src15_channel -> crosser_009:in_channel
	wire          cmd_xbar_demux_001_src15_ready;                                                                           // crosser_009:in_ready -> cmd_xbar_demux_001:src15_ready
	wire          crosser_010_out_endofpacket;                                                                              // crosser_010:out_endofpacket -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_010_out_valid;                                                                                    // crosser_010:out_valid -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_010_out_startofpacket;                                                                            // crosser_010:out_startofpacket -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_010_out_data;                                                                                     // crosser_010:out_data -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_010_out_channel;                                                                                  // crosser_010:out_channel -> baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                                     // cmd_xbar_demux_001:src16_endofpacket -> crosser_010:in_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                           // cmd_xbar_demux_001:src16_valid -> crosser_010:in_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                                   // cmd_xbar_demux_001:src16_startofpacket -> crosser_010:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src16_data;                                                                            // cmd_xbar_demux_001:src16_data -> crosser_010:in_data
	wire   [22:0] cmd_xbar_demux_001_src16_channel;                                                                         // cmd_xbar_demux_001:src16_channel -> crosser_010:in_channel
	wire          cmd_xbar_demux_001_src16_ready;                                                                           // crosser_010:in_ready -> cmd_xbar_demux_001:src16_ready
	wire          crosser_011_out_endofpacket;                                                                              // crosser_011:out_endofpacket -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_011_out_valid;                                                                                    // crosser_011:out_valid -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_011_out_startofpacket;                                                                            // crosser_011:out_startofpacket -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_011_out_data;                                                                                     // crosser_011:out_data -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_011_out_channel;                                                                                  // crosser_011:out_channel -> skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                                     // cmd_xbar_demux_001:src17_endofpacket -> crosser_011:in_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                           // cmd_xbar_demux_001:src17_valid -> crosser_011:in_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                                   // cmd_xbar_demux_001:src17_startofpacket -> crosser_011:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src17_data;                                                                            // cmd_xbar_demux_001:src17_data -> crosser_011:in_data
	wire   [22:0] cmd_xbar_demux_001_src17_channel;                                                                         // cmd_xbar_demux_001:src17_channel -> crosser_011:in_channel
	wire          cmd_xbar_demux_001_src17_ready;                                                                           // crosser_011:in_ready -> cmd_xbar_demux_001:src17_ready
	wire          crosser_012_out_endofpacket;                                                                              // crosser_012:out_endofpacket -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_012_out_valid;                                                                                    // crosser_012:out_valid -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_012_out_startofpacket;                                                                            // crosser_012:out_startofpacket -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_012_out_data;                                                                                     // crosser_012:out_data -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_012_out_channel;                                                                                  // crosser_012:out_channel -> knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                                     // cmd_xbar_demux_001:src18_endofpacket -> crosser_012:in_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                           // cmd_xbar_demux_001:src18_valid -> crosser_012:in_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                                   // cmd_xbar_demux_001:src18_startofpacket -> crosser_012:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src18_data;                                                                            // cmd_xbar_demux_001:src18_data -> crosser_012:in_data
	wire   [22:0] cmd_xbar_demux_001_src18_channel;                                                                         // cmd_xbar_demux_001:src18_channel -> crosser_012:in_channel
	wire          cmd_xbar_demux_001_src18_ready;                                                                           // crosser_012:in_ready -> cmd_xbar_demux_001:src18_ready
	wire          crosser_013_out_endofpacket;                                                                              // crosser_013:out_endofpacket -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_013_out_valid;                                                                                    // crosser_013:out_valid -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_013_out_startofpacket;                                                                            // crosser_013:out_startofpacket -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_013_out_data;                                                                                     // crosser_013:out_data -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_013_out_channel;                                                                                  // crosser_013:out_channel -> emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src19_endofpacket;                                                                     // cmd_xbar_demux_001:src19_endofpacket -> crosser_013:in_endofpacket
	wire          cmd_xbar_demux_001_src19_valid;                                                                           // cmd_xbar_demux_001:src19_valid -> crosser_013:in_valid
	wire          cmd_xbar_demux_001_src19_startofpacket;                                                                   // cmd_xbar_demux_001:src19_startofpacket -> crosser_013:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src19_data;                                                                            // cmd_xbar_demux_001:src19_data -> crosser_013:in_data
	wire   [22:0] cmd_xbar_demux_001_src19_channel;                                                                         // cmd_xbar_demux_001:src19_channel -> crosser_013:in_channel
	wire          cmd_xbar_demux_001_src19_ready;                                                                           // crosser_013:in_ready -> cmd_xbar_demux_001:src19_ready
	wire          crosser_014_out_endofpacket;                                                                              // crosser_014:out_endofpacket -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_014_out_valid;                                                                                    // crosser_014:out_valid -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_014_out_startofpacket;                                                                            // crosser_014:out_startofpacket -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_014_out_data;                                                                                     // crosser_014:out_data -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_014_out_channel;                                                                                  // crosser_014:out_channel -> EndTSetReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src20_endofpacket;                                                                     // cmd_xbar_demux_001:src20_endofpacket -> crosser_014:in_endofpacket
	wire          cmd_xbar_demux_001_src20_valid;                                                                           // cmd_xbar_demux_001:src20_valid -> crosser_014:in_valid
	wire          cmd_xbar_demux_001_src20_startofpacket;                                                                   // cmd_xbar_demux_001:src20_startofpacket -> crosser_014:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src20_data;                                                                            // cmd_xbar_demux_001:src20_data -> crosser_014:in_data
	wire   [22:0] cmd_xbar_demux_001_src20_channel;                                                                         // cmd_xbar_demux_001:src20_channel -> crosser_014:in_channel
	wire          cmd_xbar_demux_001_src20_ready;                                                                           // crosser_014:in_ready -> cmd_xbar_demux_001:src20_ready
	wire          crosser_015_out_endofpacket;                                                                              // crosser_015:out_endofpacket -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_015_out_valid;                                                                                    // crosser_015:out_valid -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_015_out_startofpacket;                                                                            // crosser_015:out_startofpacket -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_015_out_data;                                                                                     // crosser_015:out_data -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_015_out_channel;                                                                                  // crosser_015:out_channel -> FullReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src21_endofpacket;                                                                     // cmd_xbar_demux_001:src21_endofpacket -> crosser_015:in_endofpacket
	wire          cmd_xbar_demux_001_src21_valid;                                                                           // cmd_xbar_demux_001:src21_valid -> crosser_015:in_valid
	wire          cmd_xbar_demux_001_src21_startofpacket;                                                                   // cmd_xbar_demux_001:src21_startofpacket -> crosser_015:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src21_data;                                                                            // cmd_xbar_demux_001:src21_data -> crosser_015:in_data
	wire   [22:0] cmd_xbar_demux_001_src21_channel;                                                                         // cmd_xbar_demux_001:src21_channel -> crosser_015:in_channel
	wire          cmd_xbar_demux_001_src21_ready;                                                                           // crosser_015:in_ready -> cmd_xbar_demux_001:src21_ready
	wire          crosser_016_out_endofpacket;                                                                              // crosser_016:out_endofpacket -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_016_out_valid;                                                                                    // crosser_016:out_valid -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_016_out_startofpacket;                                                                            // crosser_016:out_startofpacket -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [102:0] crosser_016_out_data;                                                                                     // crosser_016:out_data -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [22:0] crosser_016_out_channel;                                                                                  // crosser_016:out_channel -> NTrReg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src22_endofpacket;                                                                     // cmd_xbar_demux_001:src22_endofpacket -> crosser_016:in_endofpacket
	wire          cmd_xbar_demux_001_src22_valid;                                                                           // cmd_xbar_demux_001:src22_valid -> crosser_016:in_valid
	wire          cmd_xbar_demux_001_src22_startofpacket;                                                                   // cmd_xbar_demux_001:src22_startofpacket -> crosser_016:in_startofpacket
	wire  [102:0] cmd_xbar_demux_001_src22_data;                                                                            // cmd_xbar_demux_001:src22_data -> crosser_016:in_data
	wire   [22:0] cmd_xbar_demux_001_src22_channel;                                                                         // cmd_xbar_demux_001:src22_channel -> crosser_016:in_channel
	wire          cmd_xbar_demux_001_src22_ready;                                                                           // crosser_016:in_ready -> cmd_xbar_demux_001:src22_ready
	wire          crosser_017_out_endofpacket;                                                                              // crosser_017:out_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          crosser_017_out_valid;                                                                                    // crosser_017:out_valid -> rsp_xbar_mux_001:sink4_valid
	wire          crosser_017_out_startofpacket;                                                                            // crosser_017:out_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [102:0] crosser_017_out_data;                                                                                     // crosser_017:out_data -> rsp_xbar_mux_001:sink4_data
	wire   [22:0] crosser_017_out_channel;                                                                                  // crosser_017:out_channel -> rsp_xbar_mux_001:sink4_channel
	wire          crosser_017_out_ready;                                                                                    // rsp_xbar_mux_001:sink4_ready -> crosser_017:out_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                      // rsp_xbar_demux_004:src0_endofpacket -> crosser_017:in_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                            // rsp_xbar_demux_004:src0_valid -> crosser_017:in_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                    // rsp_xbar_demux_004:src0_startofpacket -> crosser_017:in_startofpacket
	wire  [102:0] rsp_xbar_demux_004_src0_data;                                                                             // rsp_xbar_demux_004:src0_data -> crosser_017:in_data
	wire   [22:0] rsp_xbar_demux_004_src0_channel;                                                                          // rsp_xbar_demux_004:src0_channel -> crosser_017:in_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                            // crosser_017:in_ready -> rsp_xbar_demux_004:src0_ready
	wire          crosser_018_out_endofpacket;                                                                              // crosser_018:out_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          crosser_018_out_valid;                                                                                    // crosser_018:out_valid -> rsp_xbar_mux_001:sink7_valid
	wire          crosser_018_out_startofpacket;                                                                            // crosser_018:out_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [102:0] crosser_018_out_data;                                                                                     // crosser_018:out_data -> rsp_xbar_mux_001:sink7_data
	wire   [22:0] crosser_018_out_channel;                                                                                  // crosser_018:out_channel -> rsp_xbar_mux_001:sink7_channel
	wire          crosser_018_out_ready;                                                                                    // rsp_xbar_mux_001:sink7_ready -> crosser_018:out_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                      // rsp_xbar_demux_007:src0_endofpacket -> crosser_018:in_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                            // rsp_xbar_demux_007:src0_valid -> crosser_018:in_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                    // rsp_xbar_demux_007:src0_startofpacket -> crosser_018:in_startofpacket
	wire  [102:0] rsp_xbar_demux_007_src0_data;                                                                             // rsp_xbar_demux_007:src0_data -> crosser_018:in_data
	wire   [22:0] rsp_xbar_demux_007_src0_channel;                                                                          // rsp_xbar_demux_007:src0_channel -> crosser_018:in_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                            // crosser_018:in_ready -> rsp_xbar_demux_007:src0_ready
	wire          crosser_019_out_endofpacket;                                                                              // crosser_019:out_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          crosser_019_out_valid;                                                                                    // crosser_019:out_valid -> rsp_xbar_mux_001:sink8_valid
	wire          crosser_019_out_startofpacket;                                                                            // crosser_019:out_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [102:0] crosser_019_out_data;                                                                                     // crosser_019:out_data -> rsp_xbar_mux_001:sink8_data
	wire   [22:0] crosser_019_out_channel;                                                                                  // crosser_019:out_channel -> rsp_xbar_mux_001:sink8_channel
	wire          crosser_019_out_ready;                                                                                    // rsp_xbar_mux_001:sink8_ready -> crosser_019:out_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                      // rsp_xbar_demux_008:src0_endofpacket -> crosser_019:in_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                            // rsp_xbar_demux_008:src0_valid -> crosser_019:in_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                    // rsp_xbar_demux_008:src0_startofpacket -> crosser_019:in_startofpacket
	wire  [102:0] rsp_xbar_demux_008_src0_data;                                                                             // rsp_xbar_demux_008:src0_data -> crosser_019:in_data
	wire   [22:0] rsp_xbar_demux_008_src0_channel;                                                                          // rsp_xbar_demux_008:src0_channel -> crosser_019:in_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                            // crosser_019:in_ready -> rsp_xbar_demux_008:src0_ready
	wire          crosser_020_out_endofpacket;                                                                              // crosser_020:out_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          crosser_020_out_valid;                                                                                    // crosser_020:out_valid -> rsp_xbar_mux_001:sink9_valid
	wire          crosser_020_out_startofpacket;                                                                            // crosser_020:out_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [102:0] crosser_020_out_data;                                                                                     // crosser_020:out_data -> rsp_xbar_mux_001:sink9_data
	wire   [22:0] crosser_020_out_channel;                                                                                  // crosser_020:out_channel -> rsp_xbar_mux_001:sink9_channel
	wire          crosser_020_out_ready;                                                                                    // rsp_xbar_mux_001:sink9_ready -> crosser_020:out_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                      // rsp_xbar_demux_009:src0_endofpacket -> crosser_020:in_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                            // rsp_xbar_demux_009:src0_valid -> crosser_020:in_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                    // rsp_xbar_demux_009:src0_startofpacket -> crosser_020:in_startofpacket
	wire  [102:0] rsp_xbar_demux_009_src0_data;                                                                             // rsp_xbar_demux_009:src0_data -> crosser_020:in_data
	wire   [22:0] rsp_xbar_demux_009_src0_channel;                                                                          // rsp_xbar_demux_009:src0_channel -> crosser_020:in_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                            // crosser_020:in_ready -> rsp_xbar_demux_009:src0_ready
	wire          crosser_021_out_endofpacket;                                                                              // crosser_021:out_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          crosser_021_out_valid;                                                                                    // crosser_021:out_valid -> rsp_xbar_mux_001:sink10_valid
	wire          crosser_021_out_startofpacket;                                                                            // crosser_021:out_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [102:0] crosser_021_out_data;                                                                                     // crosser_021:out_data -> rsp_xbar_mux_001:sink10_data
	wire   [22:0] crosser_021_out_channel;                                                                                  // crosser_021:out_channel -> rsp_xbar_mux_001:sink10_channel
	wire          crosser_021_out_ready;                                                                                    // rsp_xbar_mux_001:sink10_ready -> crosser_021:out_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                      // rsp_xbar_demux_010:src0_endofpacket -> crosser_021:in_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                            // rsp_xbar_demux_010:src0_valid -> crosser_021:in_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                    // rsp_xbar_demux_010:src0_startofpacket -> crosser_021:in_startofpacket
	wire  [102:0] rsp_xbar_demux_010_src0_data;                                                                             // rsp_xbar_demux_010:src0_data -> crosser_021:in_data
	wire   [22:0] rsp_xbar_demux_010_src0_channel;                                                                          // rsp_xbar_demux_010:src0_channel -> crosser_021:in_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                            // crosser_021:in_ready -> rsp_xbar_demux_010:src0_ready
	wire          crosser_022_out_endofpacket;                                                                              // crosser_022:out_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          crosser_022_out_valid;                                                                                    // crosser_022:out_valid -> rsp_xbar_mux_001:sink11_valid
	wire          crosser_022_out_startofpacket;                                                                            // crosser_022:out_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [102:0] crosser_022_out_data;                                                                                     // crosser_022:out_data -> rsp_xbar_mux_001:sink11_data
	wire   [22:0] crosser_022_out_channel;                                                                                  // crosser_022:out_channel -> rsp_xbar_mux_001:sink11_channel
	wire          crosser_022_out_ready;                                                                                    // rsp_xbar_mux_001:sink11_ready -> crosser_022:out_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                      // rsp_xbar_demux_011:src0_endofpacket -> crosser_022:in_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                            // rsp_xbar_demux_011:src0_valid -> crosser_022:in_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                    // rsp_xbar_demux_011:src0_startofpacket -> crosser_022:in_startofpacket
	wire  [102:0] rsp_xbar_demux_011_src0_data;                                                                             // rsp_xbar_demux_011:src0_data -> crosser_022:in_data
	wire   [22:0] rsp_xbar_demux_011_src0_channel;                                                                          // rsp_xbar_demux_011:src0_channel -> crosser_022:in_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                            // crosser_022:in_ready -> rsp_xbar_demux_011:src0_ready
	wire          crosser_023_out_endofpacket;                                                                              // crosser_023:out_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          crosser_023_out_valid;                                                                                    // crosser_023:out_valid -> rsp_xbar_mux_001:sink12_valid
	wire          crosser_023_out_startofpacket;                                                                            // crosser_023:out_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [102:0] crosser_023_out_data;                                                                                     // crosser_023:out_data -> rsp_xbar_mux_001:sink12_data
	wire   [22:0] crosser_023_out_channel;                                                                                  // crosser_023:out_channel -> rsp_xbar_mux_001:sink12_channel
	wire          crosser_023_out_ready;                                                                                    // rsp_xbar_mux_001:sink12_ready -> crosser_023:out_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                      // rsp_xbar_demux_012:src0_endofpacket -> crosser_023:in_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                            // rsp_xbar_demux_012:src0_valid -> crosser_023:in_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                    // rsp_xbar_demux_012:src0_startofpacket -> crosser_023:in_startofpacket
	wire  [102:0] rsp_xbar_demux_012_src0_data;                                                                             // rsp_xbar_demux_012:src0_data -> crosser_023:in_data
	wire   [22:0] rsp_xbar_demux_012_src0_channel;                                                                          // rsp_xbar_demux_012:src0_channel -> crosser_023:in_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                            // crosser_023:in_ready -> rsp_xbar_demux_012:src0_ready
	wire          crosser_024_out_endofpacket;                                                                              // crosser_024:out_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          crosser_024_out_valid;                                                                                    // crosser_024:out_valid -> rsp_xbar_mux_001:sink13_valid
	wire          crosser_024_out_startofpacket;                                                                            // crosser_024:out_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [102:0] crosser_024_out_data;                                                                                     // crosser_024:out_data -> rsp_xbar_mux_001:sink13_data
	wire   [22:0] crosser_024_out_channel;                                                                                  // crosser_024:out_channel -> rsp_xbar_mux_001:sink13_channel
	wire          crosser_024_out_ready;                                                                                    // rsp_xbar_mux_001:sink13_ready -> crosser_024:out_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                      // rsp_xbar_demux_013:src0_endofpacket -> crosser_024:in_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                            // rsp_xbar_demux_013:src0_valid -> crosser_024:in_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                    // rsp_xbar_demux_013:src0_startofpacket -> crosser_024:in_startofpacket
	wire  [102:0] rsp_xbar_demux_013_src0_data;                                                                             // rsp_xbar_demux_013:src0_data -> crosser_024:in_data
	wire   [22:0] rsp_xbar_demux_013_src0_channel;                                                                          // rsp_xbar_demux_013:src0_channel -> crosser_024:in_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                            // crosser_024:in_ready -> rsp_xbar_demux_013:src0_ready
	wire          crosser_025_out_endofpacket;                                                                              // crosser_025:out_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          crosser_025_out_valid;                                                                                    // crosser_025:out_valid -> rsp_xbar_mux_001:sink14_valid
	wire          crosser_025_out_startofpacket;                                                                            // crosser_025:out_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [102:0] crosser_025_out_data;                                                                                     // crosser_025:out_data -> rsp_xbar_mux_001:sink14_data
	wire   [22:0] crosser_025_out_channel;                                                                                  // crosser_025:out_channel -> rsp_xbar_mux_001:sink14_channel
	wire          crosser_025_out_ready;                                                                                    // rsp_xbar_mux_001:sink14_ready -> crosser_025:out_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                      // rsp_xbar_demux_014:src0_endofpacket -> crosser_025:in_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                            // rsp_xbar_demux_014:src0_valid -> crosser_025:in_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                    // rsp_xbar_demux_014:src0_startofpacket -> crosser_025:in_startofpacket
	wire  [102:0] rsp_xbar_demux_014_src0_data;                                                                             // rsp_xbar_demux_014:src0_data -> crosser_025:in_data
	wire   [22:0] rsp_xbar_demux_014_src0_channel;                                                                          // rsp_xbar_demux_014:src0_channel -> crosser_025:in_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                            // crosser_025:in_ready -> rsp_xbar_demux_014:src0_ready
	wire          crosser_026_out_endofpacket;                                                                              // crosser_026:out_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          crosser_026_out_valid;                                                                                    // crosser_026:out_valid -> rsp_xbar_mux_001:sink15_valid
	wire          crosser_026_out_startofpacket;                                                                            // crosser_026:out_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [102:0] crosser_026_out_data;                                                                                     // crosser_026:out_data -> rsp_xbar_mux_001:sink15_data
	wire   [22:0] crosser_026_out_channel;                                                                                  // crosser_026:out_channel -> rsp_xbar_mux_001:sink15_channel
	wire          crosser_026_out_ready;                                                                                    // rsp_xbar_mux_001:sink15_ready -> crosser_026:out_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                      // rsp_xbar_demux_015:src0_endofpacket -> crosser_026:in_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                            // rsp_xbar_demux_015:src0_valid -> crosser_026:in_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                    // rsp_xbar_demux_015:src0_startofpacket -> crosser_026:in_startofpacket
	wire  [102:0] rsp_xbar_demux_015_src0_data;                                                                             // rsp_xbar_demux_015:src0_data -> crosser_026:in_data
	wire   [22:0] rsp_xbar_demux_015_src0_channel;                                                                          // rsp_xbar_demux_015:src0_channel -> crosser_026:in_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                            // crosser_026:in_ready -> rsp_xbar_demux_015:src0_ready
	wire          crosser_027_out_endofpacket;                                                                              // crosser_027:out_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          crosser_027_out_valid;                                                                                    // crosser_027:out_valid -> rsp_xbar_mux_001:sink16_valid
	wire          crosser_027_out_startofpacket;                                                                            // crosser_027:out_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [102:0] crosser_027_out_data;                                                                                     // crosser_027:out_data -> rsp_xbar_mux_001:sink16_data
	wire   [22:0] crosser_027_out_channel;                                                                                  // crosser_027:out_channel -> rsp_xbar_mux_001:sink16_channel
	wire          crosser_027_out_ready;                                                                                    // rsp_xbar_mux_001:sink16_ready -> crosser_027:out_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                      // rsp_xbar_demux_016:src0_endofpacket -> crosser_027:in_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                            // rsp_xbar_demux_016:src0_valid -> crosser_027:in_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                    // rsp_xbar_demux_016:src0_startofpacket -> crosser_027:in_startofpacket
	wire  [102:0] rsp_xbar_demux_016_src0_data;                                                                             // rsp_xbar_demux_016:src0_data -> crosser_027:in_data
	wire   [22:0] rsp_xbar_demux_016_src0_channel;                                                                          // rsp_xbar_demux_016:src0_channel -> crosser_027:in_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                            // crosser_027:in_ready -> rsp_xbar_demux_016:src0_ready
	wire          crosser_028_out_endofpacket;                                                                              // crosser_028:out_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          crosser_028_out_valid;                                                                                    // crosser_028:out_valid -> rsp_xbar_mux_001:sink17_valid
	wire          crosser_028_out_startofpacket;                                                                            // crosser_028:out_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [102:0] crosser_028_out_data;                                                                                     // crosser_028:out_data -> rsp_xbar_mux_001:sink17_data
	wire   [22:0] crosser_028_out_channel;                                                                                  // crosser_028:out_channel -> rsp_xbar_mux_001:sink17_channel
	wire          crosser_028_out_ready;                                                                                    // rsp_xbar_mux_001:sink17_ready -> crosser_028:out_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                      // rsp_xbar_demux_017:src0_endofpacket -> crosser_028:in_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                            // rsp_xbar_demux_017:src0_valid -> crosser_028:in_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                    // rsp_xbar_demux_017:src0_startofpacket -> crosser_028:in_startofpacket
	wire  [102:0] rsp_xbar_demux_017_src0_data;                                                                             // rsp_xbar_demux_017:src0_data -> crosser_028:in_data
	wire   [22:0] rsp_xbar_demux_017_src0_channel;                                                                          // rsp_xbar_demux_017:src0_channel -> crosser_028:in_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                            // crosser_028:in_ready -> rsp_xbar_demux_017:src0_ready
	wire          crosser_029_out_endofpacket;                                                                              // crosser_029:out_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          crosser_029_out_valid;                                                                                    // crosser_029:out_valid -> rsp_xbar_mux_001:sink18_valid
	wire          crosser_029_out_startofpacket;                                                                            // crosser_029:out_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [102:0] crosser_029_out_data;                                                                                     // crosser_029:out_data -> rsp_xbar_mux_001:sink18_data
	wire   [22:0] crosser_029_out_channel;                                                                                  // crosser_029:out_channel -> rsp_xbar_mux_001:sink18_channel
	wire          crosser_029_out_ready;                                                                                    // rsp_xbar_mux_001:sink18_ready -> crosser_029:out_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                      // rsp_xbar_demux_018:src0_endofpacket -> crosser_029:in_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                            // rsp_xbar_demux_018:src0_valid -> crosser_029:in_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                    // rsp_xbar_demux_018:src0_startofpacket -> crosser_029:in_startofpacket
	wire  [102:0] rsp_xbar_demux_018_src0_data;                                                                             // rsp_xbar_demux_018:src0_data -> crosser_029:in_data
	wire   [22:0] rsp_xbar_demux_018_src0_channel;                                                                          // rsp_xbar_demux_018:src0_channel -> crosser_029:in_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                            // crosser_029:in_ready -> rsp_xbar_demux_018:src0_ready
	wire          crosser_030_out_endofpacket;                                                                              // crosser_030:out_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire          crosser_030_out_valid;                                                                                    // crosser_030:out_valid -> rsp_xbar_mux_001:sink19_valid
	wire          crosser_030_out_startofpacket;                                                                            // crosser_030:out_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [102:0] crosser_030_out_data;                                                                                     // crosser_030:out_data -> rsp_xbar_mux_001:sink19_data
	wire   [22:0] crosser_030_out_channel;                                                                                  // crosser_030:out_channel -> rsp_xbar_mux_001:sink19_channel
	wire          crosser_030_out_ready;                                                                                    // rsp_xbar_mux_001:sink19_ready -> crosser_030:out_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                      // rsp_xbar_demux_019:src0_endofpacket -> crosser_030:in_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                            // rsp_xbar_demux_019:src0_valid -> crosser_030:in_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                                    // rsp_xbar_demux_019:src0_startofpacket -> crosser_030:in_startofpacket
	wire  [102:0] rsp_xbar_demux_019_src0_data;                                                                             // rsp_xbar_demux_019:src0_data -> crosser_030:in_data
	wire   [22:0] rsp_xbar_demux_019_src0_channel;                                                                          // rsp_xbar_demux_019:src0_channel -> crosser_030:in_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                            // crosser_030:in_ready -> rsp_xbar_demux_019:src0_ready
	wire          crosser_031_out_endofpacket;                                                                              // crosser_031:out_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire          crosser_031_out_valid;                                                                                    // crosser_031:out_valid -> rsp_xbar_mux_001:sink20_valid
	wire          crosser_031_out_startofpacket;                                                                            // crosser_031:out_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [102:0] crosser_031_out_data;                                                                                     // crosser_031:out_data -> rsp_xbar_mux_001:sink20_data
	wire   [22:0] crosser_031_out_channel;                                                                                  // crosser_031:out_channel -> rsp_xbar_mux_001:sink20_channel
	wire          crosser_031_out_ready;                                                                                    // rsp_xbar_mux_001:sink20_ready -> crosser_031:out_ready
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                      // rsp_xbar_demux_020:src0_endofpacket -> crosser_031:in_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                            // rsp_xbar_demux_020:src0_valid -> crosser_031:in_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                                    // rsp_xbar_demux_020:src0_startofpacket -> crosser_031:in_startofpacket
	wire  [102:0] rsp_xbar_demux_020_src0_data;                                                                             // rsp_xbar_demux_020:src0_data -> crosser_031:in_data
	wire   [22:0] rsp_xbar_demux_020_src0_channel;                                                                          // rsp_xbar_demux_020:src0_channel -> crosser_031:in_channel
	wire          rsp_xbar_demux_020_src0_ready;                                                                            // crosser_031:in_ready -> rsp_xbar_demux_020:src0_ready
	wire          crosser_032_out_endofpacket;                                                                              // crosser_032:out_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire          crosser_032_out_valid;                                                                                    // crosser_032:out_valid -> rsp_xbar_mux_001:sink21_valid
	wire          crosser_032_out_startofpacket;                                                                            // crosser_032:out_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [102:0] crosser_032_out_data;                                                                                     // crosser_032:out_data -> rsp_xbar_mux_001:sink21_data
	wire   [22:0] crosser_032_out_channel;                                                                                  // crosser_032:out_channel -> rsp_xbar_mux_001:sink21_channel
	wire          crosser_032_out_ready;                                                                                    // rsp_xbar_mux_001:sink21_ready -> crosser_032:out_ready
	wire          rsp_xbar_demux_021_src0_endofpacket;                                                                      // rsp_xbar_demux_021:src0_endofpacket -> crosser_032:in_endofpacket
	wire          rsp_xbar_demux_021_src0_valid;                                                                            // rsp_xbar_demux_021:src0_valid -> crosser_032:in_valid
	wire          rsp_xbar_demux_021_src0_startofpacket;                                                                    // rsp_xbar_demux_021:src0_startofpacket -> crosser_032:in_startofpacket
	wire  [102:0] rsp_xbar_demux_021_src0_data;                                                                             // rsp_xbar_demux_021:src0_data -> crosser_032:in_data
	wire   [22:0] rsp_xbar_demux_021_src0_channel;                                                                          // rsp_xbar_demux_021:src0_channel -> crosser_032:in_channel
	wire          rsp_xbar_demux_021_src0_ready;                                                                            // crosser_032:in_ready -> rsp_xbar_demux_021:src0_ready
	wire          crosser_033_out_endofpacket;                                                                              // crosser_033:out_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	wire          crosser_033_out_valid;                                                                                    // crosser_033:out_valid -> rsp_xbar_mux_001:sink22_valid
	wire          crosser_033_out_startofpacket;                                                                            // crosser_033:out_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	wire  [102:0] crosser_033_out_data;                                                                                     // crosser_033:out_data -> rsp_xbar_mux_001:sink22_data
	wire   [22:0] crosser_033_out_channel;                                                                                  // crosser_033:out_channel -> rsp_xbar_mux_001:sink22_channel
	wire          crosser_033_out_ready;                                                                                    // rsp_xbar_mux_001:sink22_ready -> crosser_033:out_ready
	wire          rsp_xbar_demux_022_src0_endofpacket;                                                                      // rsp_xbar_demux_022:src0_endofpacket -> crosser_033:in_endofpacket
	wire          rsp_xbar_demux_022_src0_valid;                                                                            // rsp_xbar_demux_022:src0_valid -> crosser_033:in_valid
	wire          rsp_xbar_demux_022_src0_startofpacket;                                                                    // rsp_xbar_demux_022:src0_startofpacket -> crosser_033:in_startofpacket
	wire  [102:0] rsp_xbar_demux_022_src0_data;                                                                             // rsp_xbar_demux_022:src0_data -> crosser_033:in_data
	wire   [22:0] rsp_xbar_demux_022_src0_channel;                                                                          // rsp_xbar_demux_022:src0_channel -> crosser_033:in_channel
	wire          rsp_xbar_demux_022_src0_ready;                                                                            // crosser_033:in_ready -> rsp_xbar_demux_022:src0_ready
	wire          crosser_034_out_endofpacket;                                                                              // crosser_034:out_endofpacket -> cmd_xbar_mux_025:sink1_endofpacket
	wire          crosser_034_out_valid;                                                                                    // crosser_034:out_valid -> cmd_xbar_mux_025:sink1_valid
	wire          crosser_034_out_startofpacket;                                                                            // crosser_034:out_startofpacket -> cmd_xbar_mux_025:sink1_startofpacket
	wire   [86:0] crosser_034_out_data;                                                                                     // crosser_034:out_data -> cmd_xbar_mux_025:sink1_data
	wire    [3:0] crosser_034_out_channel;                                                                                  // crosser_034:out_channel -> cmd_xbar_mux_025:sink1_channel
	wire          crosser_034_out_ready;                                                                                    // cmd_xbar_mux_025:sink1_ready -> crosser_034:out_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                      // cmd_xbar_demux_004:src0_endofpacket -> crosser_034:in_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                            // cmd_xbar_demux_004:src0_valid -> crosser_034:in_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                    // cmd_xbar_demux_004:src0_startofpacket -> crosser_034:in_startofpacket
	wire   [86:0] cmd_xbar_demux_004_src0_data;                                                                             // cmd_xbar_demux_004:src0_data -> crosser_034:in_data
	wire    [3:0] cmd_xbar_demux_004_src0_channel;                                                                          // cmd_xbar_demux_004:src0_channel -> crosser_034:in_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                            // crosser_034:in_ready -> cmd_xbar_demux_004:src0_ready
	wire          crosser_035_out_endofpacket;                                                                              // crosser_035:out_endofpacket -> cmd_xbar_mux_024:sink1_endofpacket
	wire          crosser_035_out_valid;                                                                                    // crosser_035:out_valid -> cmd_xbar_mux_024:sink1_valid
	wire          crosser_035_out_startofpacket;                                                                            // crosser_035:out_startofpacket -> cmd_xbar_mux_024:sink1_startofpacket
	wire   [86:0] crosser_035_out_data;                                                                                     // crosser_035:out_data -> cmd_xbar_mux_024:sink1_data
	wire    [3:0] crosser_035_out_channel;                                                                                  // crosser_035:out_channel -> cmd_xbar_mux_024:sink1_channel
	wire          crosser_035_out_ready;                                                                                    // cmd_xbar_mux_024:sink1_ready -> crosser_035:out_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                      // cmd_xbar_demux_005:src0_endofpacket -> crosser_035:in_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                            // cmd_xbar_demux_005:src0_valid -> crosser_035:in_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                                    // cmd_xbar_demux_005:src0_startofpacket -> crosser_035:in_startofpacket
	wire   [86:0] cmd_xbar_demux_005_src0_data;                                                                             // cmd_xbar_demux_005:src0_data -> crosser_035:in_data
	wire    [3:0] cmd_xbar_demux_005_src0_channel;                                                                          // cmd_xbar_demux_005:src0_channel -> crosser_035:in_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                            // crosser_035:in_ready -> cmd_xbar_demux_005:src0_ready
	wire          crosser_036_out_endofpacket;                                                                              // crosser_036:out_endofpacket -> cmd_xbar_mux_023:sink1_endofpacket
	wire          crosser_036_out_valid;                                                                                    // crosser_036:out_valid -> cmd_xbar_mux_023:sink1_valid
	wire          crosser_036_out_startofpacket;                                                                            // crosser_036:out_startofpacket -> cmd_xbar_mux_023:sink1_startofpacket
	wire   [86:0] crosser_036_out_data;                                                                                     // crosser_036:out_data -> cmd_xbar_mux_023:sink1_data
	wire    [3:0] crosser_036_out_channel;                                                                                  // crosser_036:out_channel -> cmd_xbar_mux_023:sink1_channel
	wire          crosser_036_out_ready;                                                                                    // cmd_xbar_mux_023:sink1_ready -> crosser_036:out_ready
	wire          cmd_xbar_demux_006_src0_endofpacket;                                                                      // cmd_xbar_demux_006:src0_endofpacket -> crosser_036:in_endofpacket
	wire          cmd_xbar_demux_006_src0_valid;                                                                            // cmd_xbar_demux_006:src0_valid -> crosser_036:in_valid
	wire          cmd_xbar_demux_006_src0_startofpacket;                                                                    // cmd_xbar_demux_006:src0_startofpacket -> crosser_036:in_startofpacket
	wire   [86:0] cmd_xbar_demux_006_src0_data;                                                                             // cmd_xbar_demux_006:src0_data -> crosser_036:in_data
	wire    [3:0] cmd_xbar_demux_006_src0_channel;                                                                          // cmd_xbar_demux_006:src0_channel -> crosser_036:in_channel
	wire          cmd_xbar_demux_006_src0_ready;                                                                            // crosser_036:in_ready -> cmd_xbar_demux_006:src0_ready
	wire          crosser_037_out_endofpacket;                                                                              // crosser_037:out_endofpacket -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_037_out_valid;                                                                                    // crosser_037:out_valid -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_037_out_startofpacket;                                                                            // crosser_037:out_startofpacket -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [86:0] crosser_037_out_data;                                                                                     // crosser_037:out_data -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] crosser_037_out_channel;                                                                                  // crosser_037:out_channel -> distancecore_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_023_src1_endofpacket;                                                                      // rsp_xbar_demux_023:src1_endofpacket -> crosser_037:in_endofpacket
	wire          rsp_xbar_demux_023_src1_valid;                                                                            // rsp_xbar_demux_023:src1_valid -> crosser_037:in_valid
	wire          rsp_xbar_demux_023_src1_startofpacket;                                                                    // rsp_xbar_demux_023:src1_startofpacket -> crosser_037:in_startofpacket
	wire   [86:0] rsp_xbar_demux_023_src1_data;                                                                             // rsp_xbar_demux_023:src1_data -> crosser_037:in_data
	wire    [3:0] rsp_xbar_demux_023_src1_channel;                                                                          // rsp_xbar_demux_023:src1_channel -> crosser_037:in_channel
	wire          rsp_xbar_demux_023_src1_ready;                                                                            // crosser_037:in_ready -> rsp_xbar_demux_023:src1_ready
	wire          crosser_038_out_endofpacket;                                                                              // crosser_038:out_endofpacket -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_038_out_valid;                                                                                    // crosser_038:out_valid -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_038_out_startofpacket;                                                                            // crosser_038:out_startofpacket -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [86:0] crosser_038_out_data;                                                                                     // crosser_038:out_data -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] crosser_038_out_channel;                                                                                  // crosser_038:out_channel -> distancecore_1_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_024_src1_endofpacket;                                                                      // rsp_xbar_demux_024:src1_endofpacket -> crosser_038:in_endofpacket
	wire          rsp_xbar_demux_024_src1_valid;                                                                            // rsp_xbar_demux_024:src1_valid -> crosser_038:in_valid
	wire          rsp_xbar_demux_024_src1_startofpacket;                                                                    // rsp_xbar_demux_024:src1_startofpacket -> crosser_038:in_startofpacket
	wire   [86:0] rsp_xbar_demux_024_src1_data;                                                                             // rsp_xbar_demux_024:src1_data -> crosser_038:in_data
	wire    [3:0] rsp_xbar_demux_024_src1_channel;                                                                          // rsp_xbar_demux_024:src1_channel -> crosser_038:in_channel
	wire          rsp_xbar_demux_024_src1_ready;                                                                            // crosser_038:in_ready -> rsp_xbar_demux_024:src1_ready
	wire          crosser_039_out_endofpacket;                                                                              // crosser_039:out_endofpacket -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_039_out_valid;                                                                                    // crosser_039:out_valid -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_039_out_startofpacket;                                                                            // crosser_039:out_startofpacket -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [86:0] crosser_039_out_data;                                                                                     // crosser_039:out_data -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] crosser_039_out_channel;                                                                                  // crosser_039:out_channel -> distancecore_2_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_025_src1_endofpacket;                                                                      // rsp_xbar_demux_025:src1_endofpacket -> crosser_039:in_endofpacket
	wire          rsp_xbar_demux_025_src1_valid;                                                                            // rsp_xbar_demux_025:src1_valid -> crosser_039:in_valid
	wire          rsp_xbar_demux_025_src1_startofpacket;                                                                    // rsp_xbar_demux_025:src1_startofpacket -> crosser_039:in_startofpacket
	wire   [86:0] rsp_xbar_demux_025_src1_data;                                                                             // rsp_xbar_demux_025:src1_data -> crosser_039:in_data
	wire    [3:0] rsp_xbar_demux_025_src1_channel;                                                                          // rsp_xbar_demux_025:src1_channel -> crosser_039:in_channel
	wire          rsp_xbar_demux_025_src1_ready;                                                                            // crosser_039:in_ready -> rsp_xbar_demux_025:src1_ready
	wire          crosser_040_out_endofpacket;                                                                              // crosser_040:out_endofpacket -> cache_0_s2_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_040_out_valid;                                                                                    // crosser_040:out_valid -> cache_0_s2_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_040_out_startofpacket;                                                                            // crosser_040:out_startofpacket -> cache_0_s2_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] crosser_040_out_data;                                                                                     // crosser_040:out_data -> cache_0_s2_translator_avalon_universal_slave_0_agent:cp_data
	wire          crosser_040_out_channel;                                                                                  // crosser_040:out_channel -> cache_0_s2_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src0_endofpacket;                                                                      // cmd_xbar_demux_007:src0_endofpacket -> crosser_040:in_endofpacket
	wire          cmd_xbar_demux_007_src0_valid;                                                                            // cmd_xbar_demux_007:src0_valid -> crosser_040:in_valid
	wire          cmd_xbar_demux_007_src0_startofpacket;                                                                    // cmd_xbar_demux_007:src0_startofpacket -> crosser_040:in_startofpacket
	wire   [84:0] cmd_xbar_demux_007_src0_data;                                                                             // cmd_xbar_demux_007:src0_data -> crosser_040:in_data
	wire    [0:0] cmd_xbar_demux_007_src0_channel;                                                                          // cmd_xbar_demux_007:src0_channel -> crosser_040:in_channel
	wire          cmd_xbar_demux_007_src0_ready;                                                                            // crosser_040:in_ready -> cmd_xbar_demux_007:src0_ready
	wire          crosser_041_out_endofpacket;                                                                              // crosser_041:out_endofpacket -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_041_out_valid;                                                                                    // crosser_041:out_valid -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_041_out_startofpacket;                                                                            // crosser_041:out_startofpacket -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [84:0] crosser_041_out_data;                                                                                     // crosser_041:out_data -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:rp_data
	wire          crosser_041_out_channel;                                                                                  // crosser_041:out_channel -> distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_026_src0_endofpacket;                                                                      // rsp_xbar_demux_026:src0_endofpacket -> crosser_041:in_endofpacket
	wire          rsp_xbar_demux_026_src0_valid;                                                                            // rsp_xbar_demux_026:src0_valid -> crosser_041:in_valid
	wire          rsp_xbar_demux_026_src0_startofpacket;                                                                    // rsp_xbar_demux_026:src0_startofpacket -> crosser_041:in_startofpacket
	wire   [84:0] rsp_xbar_demux_026_src0_data;                                                                             // rsp_xbar_demux_026:src0_data -> crosser_041:in_data
	wire    [0:0] rsp_xbar_demux_026_src0_channel;                                                                          // rsp_xbar_demux_026:src0_channel -> crosser_041:in_channel
	wire          rsp_xbar_demux_026_src0_ready;                                                                            // crosser_041:in_ready -> rsp_xbar_demux_026:src0_ready
	wire          crosser_042_out_endofpacket;                                                                              // crosser_042:out_endofpacket -> cache_1_s2_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_042_out_valid;                                                                                    // crosser_042:out_valid -> cache_1_s2_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_042_out_startofpacket;                                                                            // crosser_042:out_startofpacket -> cache_1_s2_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] crosser_042_out_data;                                                                                     // crosser_042:out_data -> cache_1_s2_translator_avalon_universal_slave_0_agent:cp_data
	wire          crosser_042_out_channel;                                                                                  // crosser_042:out_channel -> cache_1_s2_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src0_endofpacket;                                                                      // cmd_xbar_demux_008:src0_endofpacket -> crosser_042:in_endofpacket
	wire          cmd_xbar_demux_008_src0_valid;                                                                            // cmd_xbar_demux_008:src0_valid -> crosser_042:in_valid
	wire          cmd_xbar_demux_008_src0_startofpacket;                                                                    // cmd_xbar_demux_008:src0_startofpacket -> crosser_042:in_startofpacket
	wire   [84:0] cmd_xbar_demux_008_src0_data;                                                                             // cmd_xbar_demux_008:src0_data -> crosser_042:in_data
	wire    [0:0] cmd_xbar_demux_008_src0_channel;                                                                          // cmd_xbar_demux_008:src0_channel -> crosser_042:in_channel
	wire          cmd_xbar_demux_008_src0_ready;                                                                            // crosser_042:in_ready -> cmd_xbar_demux_008:src0_ready
	wire          crosser_043_out_endofpacket;                                                                              // crosser_043:out_endofpacket -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_043_out_valid;                                                                                    // crosser_043:out_valid -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_043_out_startofpacket;                                                                            // crosser_043:out_startofpacket -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [84:0] crosser_043_out_data;                                                                                     // crosser_043:out_data -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:rp_data
	wire          crosser_043_out_channel;                                                                                  // crosser_043:out_channel -> distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_027_src0_endofpacket;                                                                      // rsp_xbar_demux_027:src0_endofpacket -> crosser_043:in_endofpacket
	wire          rsp_xbar_demux_027_src0_valid;                                                                            // rsp_xbar_demux_027:src0_valid -> crosser_043:in_valid
	wire          rsp_xbar_demux_027_src0_startofpacket;                                                                    // rsp_xbar_demux_027:src0_startofpacket -> crosser_043:in_startofpacket
	wire   [84:0] rsp_xbar_demux_027_src0_data;                                                                             // rsp_xbar_demux_027:src0_data -> crosser_043:in_data
	wire    [0:0] rsp_xbar_demux_027_src0_channel;                                                                          // rsp_xbar_demux_027:src0_channel -> crosser_043:in_channel
	wire          rsp_xbar_demux_027_src0_ready;                                                                            // crosser_043:in_ready -> rsp_xbar_demux_027:src0_ready
	wire          crosser_044_out_endofpacket;                                                                              // crosser_044:out_endofpacket -> cache_2_s2_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_044_out_valid;                                                                                    // crosser_044:out_valid -> cache_2_s2_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_044_out_startofpacket;                                                                            // crosser_044:out_startofpacket -> cache_2_s2_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [84:0] crosser_044_out_data;                                                                                     // crosser_044:out_data -> cache_2_s2_translator_avalon_universal_slave_0_agent:cp_data
	wire          crosser_044_out_channel;                                                                                  // crosser_044:out_channel -> cache_2_s2_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_009_src0_endofpacket;                                                                      // cmd_xbar_demux_009:src0_endofpacket -> crosser_044:in_endofpacket
	wire          cmd_xbar_demux_009_src0_valid;                                                                            // cmd_xbar_demux_009:src0_valid -> crosser_044:in_valid
	wire          cmd_xbar_demux_009_src0_startofpacket;                                                                    // cmd_xbar_demux_009:src0_startofpacket -> crosser_044:in_startofpacket
	wire   [84:0] cmd_xbar_demux_009_src0_data;                                                                             // cmd_xbar_demux_009:src0_data -> crosser_044:in_data
	wire    [0:0] cmd_xbar_demux_009_src0_channel;                                                                          // cmd_xbar_demux_009:src0_channel -> crosser_044:in_channel
	wire          cmd_xbar_demux_009_src0_ready;                                                                            // crosser_044:in_ready -> cmd_xbar_demux_009:src0_ready
	wire          crosser_045_out_endofpacket;                                                                              // crosser_045:out_endofpacket -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_045_out_valid;                                                                                    // crosser_045:out_valid -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_045_out_startofpacket;                                                                            // crosser_045:out_startofpacket -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [84:0] crosser_045_out_data;                                                                                     // crosser_045:out_data -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:rp_data
	wire          crosser_045_out_channel;                                                                                  // crosser_045:out_channel -> distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_028_src0_endofpacket;                                                                      // rsp_xbar_demux_028:src0_endofpacket -> crosser_045:in_endofpacket
	wire          rsp_xbar_demux_028_src0_valid;                                                                            // rsp_xbar_demux_028:src0_valid -> crosser_045:in_valid
	wire          rsp_xbar_demux_028_src0_startofpacket;                                                                    // rsp_xbar_demux_028:src0_startofpacket -> crosser_045:in_startofpacket
	wire   [84:0] rsp_xbar_demux_028_src0_data;                                                                             // rsp_xbar_demux_028:src0_data -> crosser_045:in_data
	wire    [0:0] rsp_xbar_demux_028_src0_channel;                                                                          // rsp_xbar_demux_028:src0_channel -> crosser_045:in_channel
	wire          rsp_xbar_demux_028_src0_ready;                                                                            // crosser_045:in_ready -> rsp_xbar_demux_028:src0_ready
	wire          irq_mapper_receiver0_irq;                                                                                 // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                 // dma:dma_ctl_irq -> irq_mapper:receiver1_irq
	wire   [31:0] cpu_0_d_irq_irq;                                                                                          // irq_mapper:sender_irq -> cpu_0:d_irq

	nios_sys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c2_clk),                                               //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                                 // reset1.reset
	);

	nios_sys_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c2_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	nios_sys_pio_0 pio_0 (
		.clk        (altpll_0_c2_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (pio_0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_pio_0)                             // external_connection.export
	);

	usbFIFOCtrl usbfifoctrl_0 (
		.clk         (altpll_0_c0_clk),                                                        //          clock.clk
		.reset_n     (~rst_controller_001_reset_out_reset),                                    //          reset.reset_n
		.read        (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write       (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect  (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.byteenable  (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable), //               .byteenable
		.address     (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata    (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata   (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.FIFO_wr_n   (FIFO_wr_n_from_the_usbFIFOCtrl_0),                                       //    conduit_end.export
		.FIFO_rd_n   (FIFO_rd_n_from_the_usbFIFOCtrl_0),                                       //  conduit_end_1.export
		.FIFO_oe_n   (FIFO_oe_n_from_the_usbFIFOCtrl_0),                                       //  conduit_end_2.export
		.FIFO_pktend (FIFO_pktend_from_the_usbFIFOCtrl_0),                                     //  conduit_end_3.export
		.FIFO_add    (FIFO_add_from_the_usbFIFOCtrl_0),                                        //  conduit_end_4.export
		.FIFO_data   (FIFO_data_to_and_from_the_usbFIFOCtrl_0),                                //  conduit_end_5.export
		.FLAGB_n     (FLAGB_n_to_the_usbFIFOCtrl_0),                                           //  conduit_end_6.export
		.FLAGC_n     (FLAGC_n_to_the_usbFIFOCtrl_0),                                           //  conduit_end_7.export
		.led         (led_from_the_usbFIFOCtrl_0)                                              //  conduit_end_8.export
	);

	nios_sys_sdram_controller sdram_controller (
		.clk            (altpll_0_c2_clk),                                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                                  // reset.reset_n
		.az_addr        (sdram_controller_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_controller_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_controller_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_controller_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_controller_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram_0),                                         //  wire.export
		.zs_ba          (zs_ba_from_the_sdram_0),                                           //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram_0),                                        //      .export
		.zs_cke         (zs_cke_from_the_sdram_0),                                          //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram_0),                                         //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram_0),                                    //      .export
		.zs_dqm         (zs_dqm_from_the_sdram_0),                                          //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram_0),                                        //      .export
		.zs_we_n        (zs_we_n_from_the_sdram_0)                                          //      .export
	);

	nios_sys_cpu_0 cpu_0 (
		.clk           (altpll_0_c2_clk),                      //                       clk.clk
		.reset_n       (~rst_controller_reset_out_reset),      //                   reset_n.reset_n
		.d_address     (cpu_0_data_master_address),            //               data_master.address
		.d_byteenable  (cpu_0_data_master_byteenable),         //                          .byteenable
		.d_read        (cpu_0_data_master_read),               //                          .read
		.d_readdata    (cpu_0_data_master_readdata),           //                          .readdata
		.d_waitrequest (cpu_0_data_master_waitrequest),        //                          .waitrequest
		.d_write       (cpu_0_data_master_write),              //                          .write
		.d_writedata   (cpu_0_data_master_writedata),          //                          .writedata
		.i_address     (cpu_0_instruction_master_address),     //        instruction_master.address
		.i_read        (cpu_0_instruction_master_read),        //                          .read
		.i_readdata    (cpu_0_instruction_master_readdata),    //                          .readdata
		.i_waitrequest (cpu_0_instruction_master_waitrequest), //                          .waitrequest
		.d_irq         (cpu_0_d_irq_irq),                      //                     d_irq.irq
		.no_ci_readra  ()                                      // custom_instruction_master.readra
	);

	nios_sys_altpll_0 altpll_0 (
		.clk       (clk_0),                              //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (altpll_0_c0_clk),                    //                    c0.clk
		.c1        (altpll_0_c1_clk),                    //                    c1.clk
		.c2        (altpll_0_c2_clk),                    //                    c2.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	nios_sys_performance_counter_0 performance_counter_0 (
		.clk           (altpll_0_c2_clk),                                                                  //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                                  //         reset.reset_n
		.address       (performance_counter_0_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (performance_counter_0_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	nios_sys_dma dma (
		.clk                (altpll_0_c2_clk),                                                  //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                                  //              reset.reset_n
		.dma_ctl_address    (dma_control_port_slave_translator_avalon_anti_slave_0_address),    // control_port_slave.address
		.dma_ctl_chipselect (dma_control_port_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.dma_ctl_readdata   (dma_control_port_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.dma_ctl_write_n    (~dma_control_port_slave_translator_avalon_anti_slave_0_write),     //                   .write_n
		.dma_ctl_writedata  (dma_control_port_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver1_irq),                                         //                irq.irq
		.read_address       (dma_read_master_address),                                          //        read_master.address
		.read_chipselect    (dma_read_master_chipselect),                                       //                   .chipselect
		.read_read_n        (dma_read_master_read),                                             //                   .read_n
		.read_readdata      (dma_read_master_readdata),                                         //                   .readdata
		.read_readdatavalid (dma_read_master_readdatavalid),                                    //                   .readdatavalid
		.read_waitrequest   (dma_read_master_waitrequest),                                      //                   .waitrequest
		.write_address      (dma_write_master_address),                                         //       write_master.address
		.write_chipselect   (dma_write_master_chipselect),                                      //                   .chipselect
		.write_waitrequest  (dma_write_master_waitrequest),                                     //                   .waitrequest
		.write_write_n      (dma_write_master_write),                                           //                   .write_n
		.write_writedata    (dma_write_master_writedata),                                       //                   .writedata
		.write_byteenable   (dma_write_master_byteenable)                                       //                   .byteenable
	);

	nios_sys_cache_0 cache_0 (
		.clk         (altpll_0_c2_clk),                                      //   clk1.clk
		.address     (cache_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect  (cache_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken       (cache_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata    (cache_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write       (cache_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata   (cache_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable  (cache_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                       // reset1.reset
		.address2    (cache_0_s2_translator_avalon_anti_slave_0_address),    //     s2.address
		.chipselect2 (cache_0_s2_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken2      (cache_0_s2_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata2   (cache_0_s2_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write2      (cache_0_s2_translator_avalon_anti_slave_0_write),      //       .write
		.writedata2  (cache_0_s2_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable2 (cache_0_s2_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.clk2        (altpll_0_c2_clk),                                      //   clk2.clk
		.reset2      (rst_controller_reset_out_reset)                        // reset2.reset
	);

	distancecore distancecore_0 (
		.Clk          (altpll_1_c0_clk),                            //           clock.clk
		.reset_n      (~rst_controller_003_reset_out_reset),        //           reset.reset_n
		.chipselect   (distancecore_0_avalon_master_chipselect),    //   avalon_master.chipselect
		.read         (distancecore_0_avalon_master_read),          //                .read
		.write        (distancecore_0_avalon_master_write),         //                .write
		.address      (distancecore_0_avalon_master_address),       //                .address
		.readdata     (distancecore_0_avalon_master_readdata),      //                .readdata
		.writedata    (distancecore_0_avalon_master_writedata),     //                .writedata
		.waitrequest  (distancecore_0_avalon_master_waitrequest),   //                .waitrequest
		.NDim         (ndimreg_ndim0_export),                       //            NDim.export
		.Cl           (distancecore_0_cl_export),                   //              Cl.export
		.Go           (knnclasscore_go0_export),                    //              Go.export
		.EndComp      (distancecore_0_endcomp_export),              //         EndComp.export
		.NTr          (ntrreg_0_ntr_export),                        //             NTr.export
		.Full         (fullreg_0_full_export),                      //            Full.export
		.Empty        (distancecore_0_empty_export),                //           Empty.export
		.EndTSetIn    (endtsetreg_0_endtset_export),                //       EndTSetIn.export
		.EndTSetOut   (distancecore_0_endtsetout_export),           //      EndTSetOut.export
		.reset        (knnclasscore_distreset0_export),             //       DistReset.export
		.Drop         (knnclasscore_drop0_export),                  //            Drop.export
		.waitrequest1 (distancecore_0_avalon_master_1_waitrequest), // avalon_master_1.waitrequest
		.chipselect1  (distancecore_0_avalon_master_1_chipselect),  //                .chipselect
		.read1        (distancecore_0_avalon_master_1_read),        //                .read
		.write1       (distancecore_0_avalon_master_1_write),       //                .write
		.address1     (distancecore_0_avalon_master_1_address),     //                .address
		.readdata1    (distancecore_0_avalon_master_1_readdata),    //                .readdata
		.writedata1   (distancecore_0_avalon_master_1_writedata),   //                .writedata
		.QAddress     (baseqaddr_0_qaddress0_export),               //        QAddress.export
		.SkipAddr     (skipaddrreg_0_skipaddr0_export),             //        SkipAddr.export
		.Dist         (distancecore_0_dist_export),                 //            Dist.export
		.Overflow     (distancecore_0_overflow_export)              //        Overflow.export
	);

	NDimReg ndimreg (
		.clk        (altpll_1_c0_clk),                                                  //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                              //          reset.reset_n
		.read       (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.NDim0      (ndimreg_ndim0_export),                                             //          NDim0.export
		.NDim1      (ndimreg_ndim1_export),                                             //          NDim1.export
		.NDim2      (ndimreg_ndim2_export),                                             //          NDim2.export
		.NDim3      ()                                                                  //          NDim3.export
	);

	nios_sys_cache_1 cache_1 (
		.clk         (altpll_0_c2_clk),                                      //   clk1.clk
		.address     (cache_1_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect  (cache_1_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken       (cache_1_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata    (cache_1_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write       (cache_1_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata   (cache_1_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable  (cache_1_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                       // reset1.reset
		.address2    (cache_1_s2_translator_avalon_anti_slave_0_address),    //     s2.address
		.chipselect2 (cache_1_s2_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken2      (cache_1_s2_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata2   (cache_1_s2_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write2      (cache_1_s2_translator_avalon_anti_slave_0_write),      //       .write
		.writedata2  (cache_1_s2_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable2 (cache_1_s2_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.clk2        (altpll_0_c2_clk),                                      //   clk2.clk
		.reset2      (rst_controller_reset_out_reset)                        // reset2.reset
	);

	distancecore distancecore_1 (
		.Clk          (altpll_1_c0_clk),                            //           clock.clk
		.reset_n      (~rst_controller_003_reset_out_reset),        //           reset.reset_n
		.chipselect   (distancecore_1_avalon_master_chipselect),    //   avalon_master.chipselect
		.read         (distancecore_1_avalon_master_read),          //                .read
		.write        (distancecore_1_avalon_master_write),         //                .write
		.address      (distancecore_1_avalon_master_address),       //                .address
		.readdata     (distancecore_1_avalon_master_readdata),      //                .readdata
		.writedata    (distancecore_1_avalon_master_writedata),     //                .writedata
		.waitrequest  (distancecore_1_avalon_master_waitrequest),   //                .waitrequest
		.NDim         (ndimreg_ndim1_export),                       //            NDim.export
		.Cl           (distancecore_1_cl_export),                   //              Cl.export
		.Go           (knnclasscore_go1_export),                    //              Go.export
		.EndComp      (distancecore_1_endcomp_export),              //         EndComp.export
		.NTr          (ntrreg_1_ntr_export),                        //             NTr.export
		.Full         (fullreg_1_full_export),                      //            Full.export
		.Empty        (distancecore_1_empty_export),                //           Empty.export
		.EndTSetIn    (endtsetreg_1_endtset_export),                //       EndTSetIn.export
		.EndTSetOut   (distancecore_1_endtsetout_export),           //      EndTSetOut.export
		.reset        (knnclasscore_distreset1_export),             //       DistReset.export
		.Drop         (knnclasscore_drop1_export),                  //            Drop.export
		.waitrequest1 (distancecore_1_avalon_master_1_waitrequest), // avalon_master_1.waitrequest
		.chipselect1  (distancecore_1_avalon_master_1_chipselect),  //                .chipselect
		.read1        (distancecore_1_avalon_master_1_read),        //                .read
		.write1       (distancecore_1_avalon_master_1_write),       //                .write
		.address1     (distancecore_1_avalon_master_1_address),     //                .address
		.readdata1    (distancecore_1_avalon_master_1_readdata),    //                .readdata
		.writedata1   (distancecore_1_avalon_master_1_writedata),   //                .writedata
		.QAddress     (baseqaddr_0_qaddress1_export),               //        QAddress.export
		.SkipAddr     (skipaddrreg_0_skipaddr1_export),             //        SkipAddr.export
		.Dist         (distancecore_1_dist_export),                 //            Dist.export
		.Overflow     (distancecore_1_overflow_export)              //        Overflow.export
	);

	KnnWrapper knnclasscore (
		.Clk        (altpll_1_c0_clk),                                                       //          clock.clk
		.Reset      (~rst_controller_003_reset_out_reset),                                   //          reset.reset_n
		.Dist0      (distancecore_0_dist_export),                                            //          Dist0.export
		.Dist1      (distancecore_1_dist_export),                                            //          Dist1.export
		.EndComp0   (distancecore_0_endcomp_export),                                         //       EndComp0.export
		.EndComp1   (distancecore_1_endcomp_export),                                         //       EndComp1.export
		.Go0        (knnclasscore_go0_export),                                               //            Go0.export
		.Go1        (knnclasscore_go1_export),                                               //            Go1.export
		.Cl0        (distancecore_0_cl_export),                                              //            Cl0.export
		.Cl1        (distancecore_1_cl_export),                                              //            Cl1.export
		.EndTSet0   (distancecore_0_endtsetout_export),                                      //       EndTSet0.export
		.EndTSet1   (distancecore_1_endtsetout_export),                                      //       EndTSet1.export
		.DistReset0 (knnclasscore_distreset0_export),                                        //     DistReset0.export
		.DistReset1 (knnclasscore_distreset1_export),                                        //     DistReset1.export
		.Drop0      (knnclasscore_drop0_export),                                             //          Drop0.export
		.Drop1      (knnclasscore_drop1_export),                                             //          Drop1.export
		.read       (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.Overflow1  (distancecore_1_overflow_export),                                        //      Overflow1.export
		.Overflow0  (distancecore_0_overflow_export),                                        //      Overflow0.export
		.Overflow2  (distancecore_2_overflow_export),                                        //      Overflow2.export
		.Drop2      (knnclasscore_drop2_export),                                             //          Drop2.export
		.DistReset2 (knnclasscore_distreset2_export),                                        //     DistReset2.export
		.Go2        (knnclasscore_go2_export),                                               //            Go2.export
		.Dist2      (distancecore_2_dist_export),                                            //          Dist2.export
		.EndTSet2   (distancecore_2_endtsetout_export),                                      //       EndTSet2.export
		.Cl2        (distancecore_2_cl_export),                                              //            Cl2.export
		.EndComp2   (distancecore_2_endcomp_export)                                          //       EndComp2.export
	);

	EndTSetReg endtsetreg_0 (
		.clk        (altpll_1_c0_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                   //          reset.reset_n
		.read       (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.EndTSet    (endtsetreg_0_endtset_export)                                            //        EndTSet.export
	);

	FullReg fullreg_0 (
		.clk        (altpll_1_c0_clk),                                                    //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                //          reset.reset_n
		.read       (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.Full       (fullreg_0_full_export)                                               //           Full.export
	);

	FullReg fullreg_1 (
		.clk        (altpll_1_c0_clk),                                                    //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                //          reset.reset_n
		.read       (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.Full       (fullreg_1_full_export)                                               //           Full.export
	);

	NTrReg ntrreg_0 (
		.clk        (altpll_1_c0_clk),                                                   //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                               //          reset.reset_n
		.read       (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.NTr        (ntrreg_0_ntr_export)                                                //            NTr.export
	);

	NTrReg ntrreg_1 (
		.clk        (altpll_1_c0_clk),                                                   //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                               //          reset.reset_n
		.read       (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.NTr        (ntrreg_1_ntr_export)                                                //            NTr.export
	);

	EmptyReg emptyreg_0 (
		.clk        (altpll_1_c0_clk),                                                     //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                 //          reset.reset_n
		.read       (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.Empty      (distancecore_0_empty_export)                                          //          Empty.export
	);

	EmptyReg emptyreg_1 (
		.clk        (altpll_1_c0_clk),                                                     //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                 //          reset.reset_n
		.read       (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.Empty      (distancecore_1_empty_export)                                          //          Empty.export
	);

	EndTSetReg endtsetreg_1 (
		.clk        (altpll_1_c0_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                   //          reset.reset_n
		.read       (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.EndTSet    (endtsetreg_1_endtset_export)                                            //        EndTSet.export
	);

	BaseQAddr baseqaddr_0 (
		.clk        (altpll_1_c0_clk),                                                      //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                  //          reset.reset_n
		.read       (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.QAddress1  (baseqaddr_0_qaddress1_export),                                         //      QAddress1.export
		.QAddress2  (baseqaddr_0_qaddress2_export),                                         //      QAddress2.export
		.QAddress0  (baseqaddr_0_qaddress0_export)                                          //      QAddress0.export
	);

	SkipAddrReg skipaddrreg_0 (
		.clk        (altpll_1_c0_clk),                                                        //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                    //          reset.reset_n
		.read       (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.SkipAddr0  (skipaddrreg_0_skipaddr0_export),                                         //      SkipAddr0.export
		.SkipAddr1  (skipaddrreg_0_skipaddr1_export),                                         //      SkipAddr1.export
		.SkipAddr2  (skipaddrreg_0_skipaddr2_export)                                          //      SkipAddr2.export
	);

	nios_sys_altpll_1 altpll_1 (
		.clk       (clk_1_clk_in_clk),                   //       inclk_interface.clk
		.reset     (rst_controller_004_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (altpll_1_c0_clk),                    //                    c0.clk
		.areset    (),                                   //        areset_conduit.export
		.c2        (),                                   //            c2_conduit.export
		.c1        (),                                   //            c1_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	distancecore distancecore_2 (
		.Clk          (altpll_1_c0_clk),                            //           clock.clk
		.reset_n      (~rst_controller_003_reset_out_reset),        //           reset.reset_n
		.chipselect   (distancecore_2_avalon_master_chipselect),    //   avalon_master.chipselect
		.read         (distancecore_2_avalon_master_read),          //                .read
		.write        (distancecore_2_avalon_master_write),         //                .write
		.address      (distancecore_2_avalon_master_address),       //                .address
		.readdata     (distancecore_2_avalon_master_readdata),      //                .readdata
		.writedata    (distancecore_2_avalon_master_writedata),     //                .writedata
		.waitrequest  (distancecore_2_avalon_master_waitrequest),   //                .waitrequest
		.NDim         (ndimreg_ndim2_export),                       //            NDim.export
		.Cl           (distancecore_2_cl_export),                   //              Cl.export
		.Go           (knnclasscore_go2_export),                    //              Go.export
		.EndComp      (distancecore_2_endcomp_export),              //         EndComp.export
		.NTr          (ntrreg_2_ntr_export),                        //             NTr.export
		.Full         (fullreg_2_full_export),                      //            Full.export
		.Empty        (distancecore_2_empty_export),                //           Empty.export
		.EndTSetIn    (endtsetreg_2_endtset_export),                //       EndTSetIn.export
		.EndTSetOut   (distancecore_2_endtsetout_export),           //      EndTSetOut.export
		.reset        (knnclasscore_distreset2_export),             //       DistReset.export
		.Drop         (knnclasscore_drop2_export),                  //            Drop.export
		.waitrequest1 (distancecore_2_avalon_master_1_waitrequest), // avalon_master_1.waitrequest
		.chipselect1  (distancecore_2_avalon_master_1_chipselect),  //                .chipselect
		.read1        (distancecore_2_avalon_master_1_read),        //                .read
		.write1       (distancecore_2_avalon_master_1_write),       //                .write
		.address1     (distancecore_2_avalon_master_1_address),     //                .address
		.readdata1    (distancecore_2_avalon_master_1_readdata),    //                .readdata
		.writedata1   (distancecore_2_avalon_master_1_writedata),   //                .writedata
		.QAddress     (baseqaddr_0_qaddress2_export),               //        QAddress.export
		.SkipAddr     (skipaddrreg_0_skipaddr2_export),             //        SkipAddr.export
		.Dist         (distancecore_2_dist_export),                 //            Dist.export
		.Overflow     (distancecore_2_overflow_export)              //        Overflow.export
	);

	EmptyReg emptyreg_2 (
		.clk        (altpll_1_c0_clk),                                                     //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                 //          reset.reset_n
		.read       (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.Empty      (distancecore_2_empty_export)                                          //          Empty.export
	);

	EndTSetReg endtsetreg_2 (
		.clk        (altpll_1_c0_clk),                                                       //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                   //          reset.reset_n
		.read       (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.EndTSet    (endtsetreg_2_endtset_export)                                            //        EndTSet.export
	);

	FullReg fullreg_2 (
		.clk        (altpll_1_c0_clk),                                                    //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                //          reset.reset_n
		.read       (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.Full       (fullreg_2_full_export)                                               //           Full.export
	);

	NTrReg ntrreg_2 (
		.clk        (altpll_1_c0_clk),                                                   //          clock.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                               //          reset.reset_n
		.read       (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read),       // avalon_slave_0.read
		.write      (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write),      //               .write
		.chipselect (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect), //               .chipselect
		.address    (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address),    //               .address
		.readdata   (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),   //               .readdata
		.writedata  (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),  //               .writedata
		.NTr        (ntrreg_2_ntr_export)                                                //            NTr.export
	);

	nios_sys_cache_2 cache_2 (
		.clk         (altpll_0_c2_clk),                                      //   clk1.clk
		.address     (cache_2_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect  (cache_2_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken       (cache_2_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata    (cache_2_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write       (cache_2_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata   (cache_2_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable  (cache_2_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                       // reset1.reset
		.address2    (cache_2_s2_translator_avalon_anti_slave_0_address),    //     s2.address
		.chipselect2 (cache_2_s2_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken2      (cache_2_s2_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata2   (cache_2_s2_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write2      (cache_2_s2_translator_avalon_anti_slave_0_write),      //       .write
		.writedata2  (cache_2_s2_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable2 (cache_2_s2_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.clk2        (altpll_0_c2_clk),                                      //   clk2.clk
		.reset2      (rst_controller_reset_out_reset)                        // reset2.reset
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_0_instruction_master_translator (
		.clk                   (altpll_0_c2_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (cpu_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_0_instruction_master_read),                                               //                          .read
		.av_readdata           (cpu_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_readdatavalid      (),                                                                            //               (terminated)
		.av_write              (1'b0),                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.av_debugaccess        (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (26),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) cpu_0_data_master_translator (
		.clk                   (altpll_0_c2_clk),                                                      //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address           (cpu_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_0_data_master_read),                                               //                          .read
		.av_readdata           (cpu_0_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_0_data_master_write),                                              //                          .write
		.av_writedata          (cpu_0_data_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                 //               (terminated)
		.av_readdatavalid      (),                                                                     //               (terminated)
		.av_lock               (1'b0),                                                                 //               (terminated)
		.av_debugaccess        (1'b0),                                                                 //               (terminated)
		.uav_clken             (),                                                                     //               (terminated)
		.av_clken              (1'b1)                                                                  //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (26),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_read_master_translator (
		.clk                   (altpll_0_c2_clk),                                                    //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (dma_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (dma_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (dma_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (dma_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (dma_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (dma_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (dma_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (dma_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (dma_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (dma_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (dma_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (dma_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (dma_read_master_waitrequest),                                        //                          .waitrequest
		.av_chipselect         (dma_read_master_chipselect),                                         //                          .chipselect
		.av_read               (~dma_read_master_read),                                              //                          .read
		.av_readdata           (dma_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (dma_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_write              (1'b0),                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                               //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                   (altpll_0_c2_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                               //              (terminated)
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_control_port_slave_translator (
		.clk                   (altpll_0_c2_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (dma_control_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (dma_control_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (dma_control_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (dma_control_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (dma_control_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                                  //              (terminated)
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (altpll_0_c2_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_0_s1_translator (
		.clk                   (altpll_0_c2_clk),                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                    //              (terminated)
		.av_begintransfer      (),                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                    //              (terminated)
		.av_burstcount         (),                                                                    //              (terminated)
		.av_byteenable         (),                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                //              (terminated)
		.av_writebyteenable    (),                                                                    //              (terminated)
		.av_lock               (),                                                                    //              (terminated)
		.av_clken              (),                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                //              (terminated)
		.av_debugaccess        (),                                                                    //              (terminated)
		.av_outputenable       ()                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) usbfifoctrl_0_avalon_slave_0_translator (
		.clk                   (altpll_0_c0_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (usbfifoctrl_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_debugaccess        (),                                                                                        //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (23),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_controller_s1_translator (
		.clk                   (altpll_0_c2_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_controller_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_controller_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_controller_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_controller_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_controller_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_controller_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_controller_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_controller_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_controller_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                               //              (terminated)
		.av_burstcount         (),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                               //              (terminated)
		.av_lock               (),                                                                               //              (terminated)
		.av_clken              (),                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                           //              (terminated)
		.av_debugaccess        (),                                                                               //              (terminated)
		.av_outputenable       ()                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) performance_counter_0_control_slave_translator (
		.clk                   (altpll_0_c2_clk),                                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                                 //                    reset.reset
		.uav_address           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (performance_counter_0_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (performance_counter_0_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (performance_counter_0_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (performance_counter_0_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (performance_counter_0_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read               (),                                                                                               //              (terminated)
		.av_beginbursttransfer (),                                                                                               //              (terminated)
		.av_burstcount         (),                                                                                               //              (terminated)
		.av_byteenable         (),                                                                                               //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                           //              (terminated)
		.av_waitrequest        (1'b0),                                                                                           //              (terminated)
		.av_writebyteenable    (),                                                                                               //              (terminated)
		.av_lock               (),                                                                                               //              (terminated)
		.av_chipselect         (),                                                                                               //              (terminated)
		.av_clken              (),                                                                                               //              (terminated)
		.uav_clken             (1'b0),                                                                                           //              (terminated)
		.av_debugaccess        (),                                                                                               //              (terminated)
		.av_outputenable       ()                                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ndimreg_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                //                    reset.reset
		.uav_address           (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ndimreg_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                  //              (terminated)
		.av_beginbursttransfer (),                                                                                  //              (terminated)
		.av_burstcount         (),                                                                                  //              (terminated)
		.av_byteenable         (),                                                                                  //              (terminated)
		.av_readdatavalid      (1'b0),                                                                              //              (terminated)
		.av_waitrequest        (1'b0),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                                  //              (terminated)
		.av_lock               (),                                                                                  //              (terminated)
		.av_clken              (),                                                                                  //              (terminated)
		.uav_clken             (1'b0),                                                                              //              (terminated)
		.av_debugaccess        (),                                                                                  //              (terminated)
		.av_outputenable       ()                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) endtsetreg_0_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (endtsetreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fullreg_0_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (fullreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fullreg_1_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (fullreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ntrreg_0_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ntrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ntrreg_1_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ntrreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) emptyreg_0_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (emptyreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) emptyreg_1_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (emptyreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) endtsetreg_1_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (endtsetreg_1_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) baseqaddr_0_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (baseqaddr_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) skipaddrreg_0_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                         //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (skipaddrreg_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_byteenable         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_debugaccess        (),                                                                                        //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) knnclasscore_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (knnclasscore_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) emptyreg_2_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                   //                    reset.reset
		.uav_address           (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (emptyreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_byteenable         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_clken              (),                                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                                 //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) endtsetreg_2_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                        //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (endtsetreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fullreg_2_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                  //                    reset.reset
		.uav_address           (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (fullreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (26),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ntrreg_2_avalon_slave_0_translator (
		.clk                   (altpll_1_c0_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                 //                    reset.reset
		.uav_address           (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (ntrreg_2_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (13),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_write_master_translator (
		.clk                   (altpll_0_c2_clk),                                                     //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                      //                     reset.reset
		.uav_address           (dma_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (dma_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (dma_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (dma_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (dma_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (dma_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (dma_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (dma_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (dma_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (dma_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (dma_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (dma_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (dma_write_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (dma_write_master_byteenable),                                         //                          .byteenable
		.av_chipselect         (dma_write_master_chipselect),                                         //                          .chipselect
		.av_write              (~dma_write_master_write),                                             //                          .write
		.av_writedata          (dma_write_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                //               (terminated)
		.av_begintransfer      (1'b0),                                                                //               (terminated)
		.av_read               (1'b0),                                                                //               (terminated)
		.av_readdata           (),                                                                    //               (terminated)
		.av_readdatavalid      (),                                                                    //               (terminated)
		.av_lock               (1'b0),                                                                //               (terminated)
		.av_debugaccess        (1'b0),                                                                //               (terminated)
		.uav_clken             (),                                                                    //               (terminated)
		.av_clken              (1'b1)                                                                 //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) distancecore_2_avalon_master_translator (
		.clk                   (altpll_1_c0_clk),                                                                 //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                              //                     reset.reset
		.uav_address           (distancecore_2_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (distancecore_2_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (distancecore_2_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (distancecore_2_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (distancecore_2_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (distancecore_2_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (distancecore_2_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (distancecore_2_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (distancecore_2_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (distancecore_2_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (distancecore_2_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (distancecore_2_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (distancecore_2_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_chipselect         (distancecore_2_avalon_master_chipselect),                                         //                          .chipselect
		.av_read               (distancecore_2_avalon_master_read),                                               //                          .read
		.av_readdata           (distancecore_2_avalon_master_readdata),                                           //                          .readdata
		.av_write              (distancecore_2_avalon_master_write),                                              //                          .write
		.av_writedata          (distancecore_2_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                            //               (terminated)
		.av_byteenable         (4'b1111),                                                                         //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                            //               (terminated)
		.av_begintransfer      (1'b0),                                                                            //               (terminated)
		.av_readdatavalid      (),                                                                                //               (terminated)
		.av_lock               (1'b0),                                                                            //               (terminated)
		.av_debugaccess        (1'b0),                                                                            //               (terminated)
		.uav_clken             (),                                                                                //               (terminated)
		.av_clken              (1'b1)                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) distancecore_1_avalon_master_translator (
		.clk                   (altpll_1_c0_clk),                                                                 //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                              //                     reset.reset
		.uav_address           (distancecore_1_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (distancecore_1_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (distancecore_1_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (distancecore_1_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (distancecore_1_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (distancecore_1_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (distancecore_1_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (distancecore_1_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (distancecore_1_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (distancecore_1_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (distancecore_1_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (distancecore_1_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (distancecore_1_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_chipselect         (distancecore_1_avalon_master_chipselect),                                         //                          .chipselect
		.av_read               (distancecore_1_avalon_master_read),                                               //                          .read
		.av_readdata           (distancecore_1_avalon_master_readdata),                                           //                          .readdata
		.av_write              (distancecore_1_avalon_master_write),                                              //                          .write
		.av_writedata          (distancecore_1_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                            //               (terminated)
		.av_byteenable         (4'b1111),                                                                         //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                            //               (terminated)
		.av_begintransfer      (1'b0),                                                                            //               (terminated)
		.av_readdatavalid      (),                                                                                //               (terminated)
		.av_lock               (1'b0),                                                                            //               (terminated)
		.av_debugaccess        (1'b0),                                                                            //               (terminated)
		.uav_clken             (),                                                                                //               (terminated)
		.av_clken              (1'b1)                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) distancecore_0_avalon_master_translator (
		.clk                   (altpll_1_c0_clk),                                                                 //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                              //                     reset.reset
		.uav_address           (distancecore_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (distancecore_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (distancecore_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (distancecore_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (distancecore_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (distancecore_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (distancecore_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (distancecore_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (distancecore_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (distancecore_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (distancecore_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (distancecore_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (distancecore_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_chipselect         (distancecore_0_avalon_master_chipselect),                                         //                          .chipselect
		.av_read               (distancecore_0_avalon_master_read),                                               //                          .read
		.av_readdata           (distancecore_0_avalon_master_readdata),                                           //                          .readdata
		.av_write              (distancecore_0_avalon_master_write),                                              //                          .write
		.av_writedata          (distancecore_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                            //               (terminated)
		.av_byteenable         (4'b1111),                                                                         //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                            //               (terminated)
		.av_begintransfer      (1'b0),                                                                            //               (terminated)
		.av_readdatavalid      (),                                                                                //               (terminated)
		.av_lock               (1'b0),                                                                            //               (terminated)
		.av_debugaccess        (1'b0),                                                                            //               (terminated)
		.uav_clken             (),                                                                                //               (terminated)
		.av_clken              (1'b1)                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cache_0_s1_translator (
		.clk                   (altpll_0_c2_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cache_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cache_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cache_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cache_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (cache_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cache_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (cache_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cache_1_s1_translator (
		.clk                   (altpll_0_c2_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cache_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cache_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cache_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cache_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (cache_1_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cache_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (cache_1_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cache_2_s1_translator (
		.clk                   (altpll_0_c2_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cache_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cache_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cache_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cache_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (cache_2_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cache_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (cache_2_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) distancecore_0_avalon_master_1_translator (
		.clk                   (altpll_1_c0_clk),                                                                   //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                //                     reset.reset
		.uav_address           (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (distancecore_0_avalon_master_1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (distancecore_0_avalon_master_1_waitrequest),                                        //                          .waitrequest
		.av_chipselect         (distancecore_0_avalon_master_1_chipselect),                                         //                          .chipselect
		.av_read               (distancecore_0_avalon_master_1_read),                                               //                          .read
		.av_readdata           (distancecore_0_avalon_master_1_readdata),                                           //                          .readdata
		.av_write              (distancecore_0_avalon_master_1_write),                                              //                          .write
		.av_writedata          (distancecore_0_avalon_master_1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                              //               (terminated)
		.av_byteenable         (4'b1111),                                                                           //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                              //               (terminated)
		.av_begintransfer      (1'b0),                                                                              //               (terminated)
		.av_readdatavalid      (),                                                                                  //               (terminated)
		.av_lock               (1'b0),                                                                              //               (terminated)
		.av_debugaccess        (1'b0),                                                                              //               (terminated)
		.uav_clken             (),                                                                                  //               (terminated)
		.av_clken              (1'b1)                                                                               //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cache_0_s2_translator (
		.clk                   (altpll_0_c2_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cache_0_s2_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cache_0_s2_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cache_0_s2_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cache_0_s2_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (cache_0_s2_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cache_0_s2_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (cache_0_s2_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) distancecore_1_avalon_master_1_translator (
		.clk                   (altpll_1_c0_clk),                                                                   //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                //                     reset.reset
		.uav_address           (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (distancecore_1_avalon_master_1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (distancecore_1_avalon_master_1_waitrequest),                                        //                          .waitrequest
		.av_chipselect         (distancecore_1_avalon_master_1_chipselect),                                         //                          .chipselect
		.av_read               (distancecore_1_avalon_master_1_read),                                               //                          .read
		.av_readdata           (distancecore_1_avalon_master_1_readdata),                                           //                          .readdata
		.av_write              (distancecore_1_avalon_master_1_write),                                              //                          .write
		.av_writedata          (distancecore_1_avalon_master_1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                              //               (terminated)
		.av_byteenable         (4'b1111),                                                                           //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                              //               (terminated)
		.av_begintransfer      (1'b0),                                                                              //               (terminated)
		.av_readdatavalid      (),                                                                                  //               (terminated)
		.av_lock               (1'b0),                                                                              //               (terminated)
		.av_debugaccess        (1'b0),                                                                              //               (terminated)
		.uav_clken             (),                                                                                  //               (terminated)
		.av_clken              (1'b1)                                                                               //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cache_1_s2_translator (
		.clk                   (altpll_0_c2_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cache_1_s2_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cache_1_s2_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cache_1_s2_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cache_1_s2_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (cache_1_s2_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cache_1_s2_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (cache_1_s2_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) distancecore_2_avalon_master_1_translator (
		.clk                   (altpll_1_c0_clk),                                                                   //                       clk.clk
		.reset                 (rst_controller_003_reset_out_reset),                                                //                     reset.reset
		.uav_address           (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (distancecore_2_avalon_master_1_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (distancecore_2_avalon_master_1_waitrequest),                                        //                          .waitrequest
		.av_chipselect         (distancecore_2_avalon_master_1_chipselect),                                         //                          .chipselect
		.av_read               (distancecore_2_avalon_master_1_read),                                               //                          .read
		.av_readdata           (distancecore_2_avalon_master_1_readdata),                                           //                          .readdata
		.av_write              (distancecore_2_avalon_master_1_write),                                              //                          .write
		.av_writedata          (distancecore_2_avalon_master_1_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                              //               (terminated)
		.av_byteenable         (4'b1111),                                                                           //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                              //               (terminated)
		.av_begintransfer      (1'b0),                                                                              //               (terminated)
		.av_readdatavalid      (),                                                                                  //               (terminated)
		.av_lock               (1'b0),                                                                              //               (terminated)
		.av_debugaccess        (1'b0),                                                                              //               (terminated)
		.uav_clken             (),                                                                                  //               (terminated)
		.av_clken              (1'b1)                                                                               //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cache_2_s2_translator (
		.clk                   (altpll_0_c2_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (cache_2_s2_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (cache_2_s2_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (cache_2_s2_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (cache_2_s2_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (cache_2_s2_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (cache_2_s2_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (cache_2_s2_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (23),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) cpu_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c2_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (cpu_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_src_valid),                                                               //        rp.valid
		.rp_data          (rsp_xbar_mux_src_data),                                                                //          .data
		.rp_channel       (rsp_xbar_mux_src_channel),                                                             //          .channel
		.rp_startofpacket (rsp_xbar_mux_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_src_endofpacket),                                                         //          .endofpacket
		.rp_ready         (rsp_xbar_mux_src_ready)                                                                //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (23),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c2_clk),                                                               //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address       (cpu_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                    //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                     //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                  //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                              //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_BEGIN_BURST           (81),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.PKT_BURST_TYPE_H          (78),
		.PKT_BURST_TYPE_L          (77),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_TRANS_EXCLUSIVE       (67),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_THREAD_ID_H           (93),
		.PKT_THREAD_ID_L           (93),
		.PKT_CACHE_H               (100),
		.PKT_CACHE_L               (97),
		.PKT_DATA_SIDEBAND_H       (80),
		.PKT_DATA_SIDEBAND_L       (80),
		.PKT_QOS_H                 (82),
		.PKT_QOS_L                 (82),
		.PKT_ADDR_SIDEBAND_H       (79),
		.PKT_ADDR_SIDEBAND_L       (79),
		.ST_DATA_W                 (103),
		.ST_CHANNEL_W              (23),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) dma_read_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c2_clk),                                                             //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address       (dma_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (dma_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (dma_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (dma_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (dma_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (dma_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (dma_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (dma_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (dma_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (dma_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (dma_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_005_src1_valid),                                               //        rp.valid
		.rp_data          (rsp_xbar_demux_005_src1_data),                                                //          .data
		.rp_channel       (rsp_xbar_demux_005_src1_channel),                                             //          .channel
		.rp_startofpacket (rsp_xbar_demux_005_src1_startofpacket),                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),                                         //          .endofpacket
		.rp_ready         (rsp_xbar_demux_005_src1_ready)                                                //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                 //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) dma_control_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                                //                .channel
		.rf_sink_ready           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                               //                .channel
		.rf_sink_ready           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (43),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (44),
		.PKT_TRANS_POSTED          (45),
		.PKT_TRANS_WRITE           (46),
		.PKT_TRANS_READ            (47),
		.PKT_TRANS_LOCK            (48),
		.PKT_SRC_ID_H              (69),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (70),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (50),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (16),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                                        // (terminated)
		.out_startofpacket (),                                                                                            // (terminated)
		.out_endofpacket   (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_controller_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                             //                .channel
		.rf_sink_ready           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (7),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                           //       clk_reset.reset
		.m0_address              (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                                          //                .channel
		.rf_sink_ready           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                           // clk_reset.reset
		.in_data           (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                                     // (terminated)
		.csr_readdata      (),                                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                     // (terminated)
		.almost_full_data  (),                                                                                                         // (terminated)
		.almost_empty_data (),                                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                                     // (terminated)
		.out_empty         (),                                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                                     // (terminated)
		.out_error         (),                                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                                     // (terminated)
		.out_channel       ()                                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_001_out_ready),                                                                       //              cp.ready
		.cp_valid                (crosser_001_out_valid),                                                                       //                .valid
		.cp_data                 (crosser_001_out_data),                                                                        //                .data
		.cp_startofpacket        (crosser_001_out_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (crosser_001_out_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (crosser_001_out_channel),                                                                     //                .channel
		.rf_sink_ready           (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                             //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                       //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_startofpacket  (1'b0),                                                                                  // (terminated)
		.in_endofpacket    (1'b0),                                                                                  // (terminated)
		.out_startofpacket (),                                                                                      // (terminated)
		.out_endofpacket   (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_002_out_ready),                                                                            //              cp.ready
		.cp_valid                (crosser_002_out_valid),                                                                            //                .valid
		.cp_data                 (crosser_002_out_data),                                                                             //                .data
		.cp_startofpacket        (crosser_002_out_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (crosser_002_out_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (crosser_002_out_channel),                                                                          //                .channel
		.rf_sink_ready           (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_003_out_ready),                                                                         //              cp.ready
		.cp_valid                (crosser_003_out_valid),                                                                         //                .valid
		.cp_data                 (crosser_003_out_data),                                                                          //                .data
		.cp_startofpacket        (crosser_003_out_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (crosser_003_out_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (crosser_003_out_channel),                                                                       //                .channel
		.rf_sink_ready           (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                               //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_004_out_ready),                                                                         //              cp.ready
		.cp_valid                (crosser_004_out_valid),                                                                         //                .valid
		.cp_data                 (crosser_004_out_data),                                                                          //                .data
		.cp_startofpacket        (crosser_004_out_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (crosser_004_out_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (crosser_004_out_channel),                                                                       //                .channel
		.rf_sink_ready           (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                               //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_005_out_ready),                                                                        //              cp.ready
		.cp_valid                (crosser_005_out_valid),                                                                        //                .valid
		.cp_data                 (crosser_005_out_data),                                                                         //                .data
		.cp_startofpacket        (crosser_005_out_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (crosser_005_out_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (crosser_005_out_channel),                                                                      //                .channel
		.rf_sink_ready           (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_startofpacket  (1'b0),                                                                                   // (terminated)
		.in_endofpacket    (1'b0),                                                                                   // (terminated)
		.out_startofpacket (),                                                                                       // (terminated)
		.out_endofpacket   (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_006_out_ready),                                                                        //              cp.ready
		.cp_valid                (crosser_006_out_valid),                                                                        //                .valid
		.cp_data                 (crosser_006_out_data),                                                                         //                .data
		.cp_startofpacket        (crosser_006_out_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (crosser_006_out_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (crosser_006_out_channel),                                                                      //                .channel
		.rf_sink_ready           (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_startofpacket  (1'b0),                                                                                   // (terminated)
		.in_endofpacket    (1'b0),                                                                                   // (terminated)
		.out_startofpacket (),                                                                                       // (terminated)
		.out_endofpacket   (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_007_out_ready),                                                                          //              cp.ready
		.cp_valid                (crosser_007_out_valid),                                                                          //                .valid
		.cp_data                 (crosser_007_out_data),                                                                           //                .data
		.cp_startofpacket        (crosser_007_out_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (crosser_007_out_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (crosser_007_out_channel),                                                                        //                .channel
		.rf_sink_ready           (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                                     // (terminated)
		.out_startofpacket (),                                                                                         // (terminated)
		.out_endofpacket   (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_008_out_ready),                                                                          //              cp.ready
		.cp_valid                (crosser_008_out_valid),                                                                          //                .valid
		.cp_data                 (crosser_008_out_data),                                                                           //                .data
		.cp_startofpacket        (crosser_008_out_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (crosser_008_out_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (crosser_008_out_channel),                                                                        //                .channel
		.rf_sink_ready           (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                                     // (terminated)
		.out_startofpacket (),                                                                                         // (terminated)
		.out_endofpacket   (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_009_out_ready),                                                                            //              cp.ready
		.cp_valid                (crosser_009_out_valid),                                                                            //                .valid
		.cp_data                 (crosser_009_out_data),                                                                             //                .data
		.cp_startofpacket        (crosser_009_out_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (crosser_009_out_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (crosser_009_out_channel),                                                                          //                .channel
		.rf_sink_ready           (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_010_out_ready),                                                                           //              cp.ready
		.cp_valid                (crosser_010_out_valid),                                                                           //                .valid
		.cp_data                 (crosser_010_out_data),                                                                            //                .data
		.cp_startofpacket        (crosser_010_out_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (crosser_010_out_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (crosser_010_out_channel),                                                                         //                .channel
		.rf_sink_ready           (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                           //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                                      // (terminated)
		.out_startofpacket (),                                                                                          // (terminated)
		.out_endofpacket   (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                   //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_011_out_ready),                                                                             //              cp.ready
		.cp_valid                (crosser_011_out_valid),                                                                             //                .valid
		.cp_data                 (crosser_011_out_data),                                                                              //                .data
		.cp_startofpacket        (crosser_011_out_startofpacket),                                                                     //                .startofpacket
		.cp_endofpacket          (crosser_011_out_endofpacket),                                                                       //                .endofpacket
		.cp_channel              (crosser_011_out_channel),                                                                           //                .channel
		.rf_sink_ready           (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                   //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                             //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                       // (terminated)
		.csr_read          (1'b0),                                                                                        // (terminated)
		.csr_write         (1'b0),                                                                                        // (terminated)
		.csr_readdata      (),                                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                        // (terminated)
		.almost_full_data  (),                                                                                            // (terminated)
		.almost_empty_data (),                                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                                        // (terminated)
		.out_startofpacket (),                                                                                            // (terminated)
		.out_endofpacket   (),                                                                                            // (terminated)
		.in_empty          (1'b0),                                                                                        // (terminated)
		.out_empty         (),                                                                                            // (terminated)
		.in_error          (1'b0),                                                                                        // (terminated)
		.out_error         (),                                                                                            // (terminated)
		.in_channel        (1'b0),                                                                                        // (terminated)
		.out_channel       ()                                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_012_out_ready),                                                                            //              cp.ready
		.cp_valid                (crosser_012_out_valid),                                                                            //                .valid
		.cp_data                 (crosser_012_out_data),                                                                             //                .data
		.cp_startofpacket        (crosser_012_out_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (crosser_012_out_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (crosser_012_out_channel),                                                                          //                .channel
		.rf_sink_ready           (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_013_out_ready),                                                                          //              cp.ready
		.cp_valid                (crosser_013_out_valid),                                                                          //                .valid
		.cp_data                 (crosser_013_out_data),                                                                           //                .data
		.cp_startofpacket        (crosser_013_out_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (crosser_013_out_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (crosser_013_out_channel),                                                                        //                .channel
		.rf_sink_ready           (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                                     // (terminated)
		.out_startofpacket (),                                                                                         // (terminated)
		.out_endofpacket   (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_014_out_ready),                                                                            //              cp.ready
		.cp_valid                (crosser_014_out_valid),                                                                            //                .valid
		.cp_data                 (crosser_014_out_data),                                                                             //                .data
		.cp_startofpacket        (crosser_014_out_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (crosser_014_out_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (crosser_014_out_channel),                                                                          //                .channel
		.rf_sink_ready           (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_015_out_ready),                                                                         //              cp.ready
		.cp_valid                (crosser_015_out_valid),                                                                         //                .valid
		.cp_data                 (crosser_015_out_data),                                                                          //                .data
		.cp_startofpacket        (crosser_015_out_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (crosser_015_out_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (crosser_015_out_channel),                                                                       //                .channel
		.rf_sink_ready           (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                               //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (81),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (61),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (62),
		.PKT_TRANS_POSTED          (63),
		.PKT_TRANS_WRITE           (64),
		.PKT_TRANS_READ            (65),
		.PKT_TRANS_LOCK            (66),
		.PKT_SRC_ID_H              (87),
		.PKT_SRC_ID_L              (83),
		.PKT_DEST_ID_H             (92),
		.PKT_DEST_ID_L             (88),
		.PKT_BURSTWRAP_H           (73),
		.PKT_BURSTWRAP_L           (71),
		.PKT_BYTE_CNT_H            (70),
		.PKT_BYTE_CNT_L            (68),
		.PKT_PROTECTION_H          (96),
		.PKT_PROTECTION_L          (94),
		.PKT_RESPONSE_STATUS_H     (102),
		.PKT_RESPONSE_STATUS_L     (101),
		.PKT_BURST_SIZE_H          (76),
		.PKT_BURST_SIZE_L          (74),
		.ST_CHANNEL_W              (23),
		.ST_DATA_W                 (103),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_1_c0_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_016_out_ready),                                                                        //              cp.ready
		.cp_valid                (crosser_016_out_valid),                                                                        //                .valid
		.cp_data                 (crosser_016_out_data),                                                                         //                .data
		.cp_startofpacket        (crosser_016_out_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (crosser_016_out_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (crosser_016_out_channel),                                                                      //                .channel
		.rf_sink_ready           (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (104),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_1_c0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_1_c0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_startofpacket  (1'b0),                                                                                   // (terminated)
		.in_endofpacket    (1'b0),                                                                                   // (terminated)
		.out_startofpacket (),                                                                                       // (terminated)
		.out_endofpacket   (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (75),
		.PKT_THREAD_ID_H           (77),
		.PKT_THREAD_ID_L           (77),
		.PKT_CACHE_H               (84),
		.PKT_CACHE_L               (81),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) dma_write_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c2_clk),                                                              //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.av_address       (dma_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (dma_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (dma_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (dma_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (dma_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (dma_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (dma_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (dma_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (dma_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (dma_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (dma_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_003_src_valid),                                                   //        rp.valid
		.rp_data          (rsp_xbar_mux_003_src_data),                                                    //          .data
		.rp_channel       (rsp_xbar_mux_003_src_channel),                                                 //          .channel
		.rp_startofpacket (rsp_xbar_mux_003_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_003_src_endofpacket),                                             //          .endofpacket
		.rp_ready         (rsp_xbar_mux_003_src_ready)                                                    //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (75),
		.PKT_THREAD_ID_H           (77),
		.PKT_THREAD_ID_L           (77),
		.PKT_CACHE_H               (84),
		.PKT_CACHE_L               (81),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) distancecore_2_avalon_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (distancecore_2_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (distancecore_2_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (distancecore_2_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (distancecore_2_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (distancecore_2_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (distancecore_2_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (distancecore_2_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (distancecore_2_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (distancecore_2_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (distancecore_2_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (distancecore_2_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (crosser_039_out_valid),                                                                    //        rp.valid
		.rp_data          (crosser_039_out_data),                                                                     //          .data
		.rp_channel       (crosser_039_out_channel),                                                                  //          .channel
		.rp_startofpacket (crosser_039_out_startofpacket),                                                            //          .startofpacket
		.rp_endofpacket   (crosser_039_out_endofpacket),                                                              //          .endofpacket
		.rp_ready         (crosser_039_out_ready)                                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (75),
		.PKT_THREAD_ID_H           (77),
		.PKT_THREAD_ID_L           (77),
		.PKT_CACHE_H               (84),
		.PKT_CACHE_L               (81),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) distancecore_1_avalon_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (distancecore_1_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (distancecore_1_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (distancecore_1_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (distancecore_1_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (distancecore_1_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (distancecore_1_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (distancecore_1_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (distancecore_1_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (distancecore_1_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (distancecore_1_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (distancecore_1_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (crosser_038_out_valid),                                                                    //        rp.valid
		.rp_data          (crosser_038_out_data),                                                                     //          .data
		.rp_channel       (crosser_038_out_channel),                                                                  //          .channel
		.rp_startofpacket (crosser_038_out_startofpacket),                                                            //          .startofpacket
		.rp_endofpacket   (crosser_038_out_endofpacket),                                                              //          .endofpacket
		.rp_ready         (crosser_038_out_ready)                                                                     //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (75),
		.PKT_THREAD_ID_H           (77),
		.PKT_THREAD_ID_L           (77),
		.PKT_CACHE_H               (84),
		.PKT_CACHE_L               (81),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (87),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) distancecore_0_avalon_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (distancecore_0_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (distancecore_0_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (distancecore_0_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (distancecore_0_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (distancecore_0_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (distancecore_0_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (distancecore_0_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (distancecore_0_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (distancecore_0_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (distancecore_0_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (distancecore_0_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (crosser_037_out_valid),                                                                    //        rp.valid
		.rp_data          (crosser_037_out_data),                                                                     //          .data
		.rp_channel       (crosser_037_out_channel),                                                                  //          .channel
		.rp_startofpacket (crosser_037_out_startofpacket),                                                            //          .startofpacket
		.rp_endofpacket   (crosser_037_out_endofpacket),                                                              //          .endofpacket
		.rp_ready         (crosser_037_out_ready)                                                                     //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_RESPONSE_STATUS_H     (86),
		.PKT_RESPONSE_STATUS_L     (85),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cache_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cache_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_023_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_023_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_023_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_023_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_023_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_023_src_channel),                                                    //                .channel
		.rf_sink_ready           (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cache_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cache_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.in_data           (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cache_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_RESPONSE_STATUS_H     (86),
		.PKT_RESPONSE_STATUS_L     (85),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cache_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cache_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_024_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_024_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_024_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_024_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_024_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_024_src_channel),                                                    //                .channel
		.rf_sink_ready           (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cache_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cache_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.in_data           (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cache_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (76),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (80),
		.PKT_PROTECTION_L          (78),
		.PKT_RESPONSE_STATUS_H     (86),
		.PKT_RESPONSE_STATUS_L     (85),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (87),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cache_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cache_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_025_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_025_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_025_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_025_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_025_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_025_src_channel),                                                    //                .channel
		.rf_sink_ready           (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (88),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cache_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cache_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.in_data           (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cache_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (74),
		.PKT_THREAD_ID_H           (75),
		.PKT_THREAD_ID_L           (75),
		.PKT_CACHE_H               (82),
		.PKT_CACHE_L               (79),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent (
		.clk              (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.av_address       (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (crosser_041_out_valid),                                                                      //        rp.valid
		.rp_data          (crosser_041_out_data),                                                                       //          .data
		.rp_channel       (crosser_041_out_channel),                                                                    //          .channel
		.rp_startofpacket (crosser_041_out_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket   (crosser_041_out_endofpacket),                                                                //          .endofpacket
		.rp_ready         (crosser_041_out_ready)                                                                       //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (74),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cache_0_s2_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cache_0_s2_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_040_out_ready),                                                           //              cp.ready
		.cp_valid                (crosser_040_out_valid),                                                           //                .valid
		.cp_data                 (crosser_040_out_data),                                                            //                .data
		.cp_startofpacket        (crosser_040_out_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (crosser_040_out_endofpacket),                                                     //                .endofpacket
		.cp_channel              (crosser_040_out_channel),                                                         //                .channel
		.rf_sink_ready           (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cache_0_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cache_0_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.in_data           (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cache_0_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (74),
		.PKT_THREAD_ID_H           (75),
		.PKT_THREAD_ID_L           (75),
		.PKT_CACHE_H               (82),
		.PKT_CACHE_L               (79),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent (
		.clk              (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.av_address       (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (crosser_043_out_valid),                                                                      //        rp.valid
		.rp_data          (crosser_043_out_data),                                                                       //          .data
		.rp_channel       (crosser_043_out_channel),                                                                    //          .channel
		.rp_startofpacket (crosser_043_out_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket   (crosser_043_out_endofpacket),                                                                //          .endofpacket
		.rp_ready         (crosser_043_out_ready)                                                                       //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (74),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cache_1_s2_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cache_1_s2_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_042_out_ready),                                                           //              cp.ready
		.cp_valid                (crosser_042_out_valid),                                                           //                .valid
		.cp_data                 (crosser_042_out_data),                                                            //                .data
		.cp_startofpacket        (crosser_042_out_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (crosser_042_out_endofpacket),                                                     //                .endofpacket
		.cp_channel              (crosser_042_out_channel),                                                         //                .channel
		.rf_sink_ready           (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cache_1_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cache_1_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.in_data           (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cache_1_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (74),
		.PKT_THREAD_ID_H           (75),
		.PKT_THREAD_ID_L           (75),
		.PKT_CACHE_H               (82),
		.PKT_CACHE_L               (79),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent (
		.clk              (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset            (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.av_address       (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (crosser_045_out_valid),                                                                      //        rp.valid
		.rp_data          (crosser_045_out_data),                                                                       //          .data
		.rp_channel       (crosser_045_out_channel),                                                                    //          .channel
		.rp_startofpacket (crosser_045_out_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket   (crosser_045_out_endofpacket),                                                                //          .endofpacket
		.rp_ready         (crosser_045_out_ready)                                                                       //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (73),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (74),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (78),
		.PKT_PROTECTION_L          (76),
		.PKT_RESPONSE_STATUS_H     (84),
		.PKT_RESPONSE_STATUS_L     (83),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (85),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) cache_2_s2_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c2_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cache_2_s2_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_044_out_ready),                                                           //              cp.ready
		.cp_valid                (crosser_044_out_valid),                                                           //                .valid
		.cp_data                 (crosser_044_out_data),                                                            //                .data
		.cp_startofpacket        (crosser_044_out_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (crosser_044_out_endofpacket),                                                     //                .endofpacket
		.cp_channel              (crosser_044_out_channel),                                                         //                .channel
		.rf_sink_ready           (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (86),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c2_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cache_2_s2_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cache_2_s2_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c2_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.in_data           (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cache_2_s2_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	nios_sys_addr_router addr_router (
		.sink_ready         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	nios_sys_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	nios_sys_addr_router_002 addr_router_002 (
		.sink_ready         (dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                   //          .valid
		.src_data           (addr_router_002_src_data),                                                    //          .data
		.src_channel        (addr_router_002_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                              //          .endofpacket
	);

	nios_sys_id_router id_router (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                            //       src.ready
		.src_valid          (id_router_src_valid),                                                            //          .valid
		.src_data           (id_router_src_data),                                                             //          .data
		.src_channel        (id_router_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                       //          .endofpacket
	);

	nios_sys_id_router id_router_001 (
		.sink_ready         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                           //       src.ready
		.src_valid          (id_router_001_src_valid),                                                           //          .valid
		.src_data           (id_router_001_src_data),                                                            //          .data
		.src_channel        (id_router_001_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                      //          .endofpacket
	);

	nios_sys_id_router_002 id_router_002 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                  //          .valid
		.src_data           (id_router_002_src_data),                                                                   //          .data
		.src_channel        (id_router_002_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                             //          .endofpacket
	);

	nios_sys_id_router_002 id_router_003 (
		.sink_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                             //          .valid
		.src_data           (id_router_003_src_data),                                              //          .data
		.src_channel        (id_router_003_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                        //          .endofpacket
	);

	nios_sys_id_router_004 id_router_004 (
		.sink_ready         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (usbfifoctrl_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                 //          .valid
		.src_data           (id_router_004_src_data),                                                                  //          .data
		.src_channel        (id_router_004_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                            //          .endofpacket
	);

	nios_sys_id_router_005 id_router_005 (
		.sink_ready         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_controller_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                        //       src.ready
		.src_valid          (id_router_005_src_valid),                                                        //          .valid
		.src_data           (id_router_005_src_data),                                                         //          .data
		.src_channel        (id_router_005_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                   //          .endofpacket
	);

	nios_sys_id_router_002 id_router_006 (
		.sink_ready         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (performance_counter_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                        //          .valid
		.src_data           (id_router_006_src_data),                                                                         //          .data
		.src_channel        (id_router_006_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                   //          .endofpacket
	);

	nios_sys_id_router_002 id_router_007 (
		.sink_ready         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ndimreg_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                   //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                           //       src.ready
		.src_valid          (id_router_007_src_valid),                                                           //          .valid
		.src_data           (id_router_007_src_data),                                                            //          .data
		.src_channel        (id_router_007_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                      //          .endofpacket
	);

	nios_sys_id_router_002 id_router_008 (
		.sink_ready         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (endtsetreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                        //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                //          .valid
		.src_data           (id_router_008_src_data),                                                                 //          .data
		.src_channel        (id_router_008_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                           //          .endofpacket
	);

	nios_sys_id_router_002 id_router_009 (
		.sink_ready         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fullreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                     //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                             //       src.ready
		.src_valid          (id_router_009_src_valid),                                                             //          .valid
		.src_data           (id_router_009_src_data),                                                              //          .data
		.src_channel        (id_router_009_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                        //          .endofpacket
	);

	nios_sys_id_router_002 id_router_010 (
		.sink_ready         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fullreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                     //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                             //       src.ready
		.src_valid          (id_router_010_src_valid),                                                             //          .valid
		.src_data           (id_router_010_src_data),                                                              //          .data
		.src_channel        (id_router_010_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                        //          .endofpacket
	);

	nios_sys_id_router_002 id_router_011 (
		.sink_ready         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ntrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                            //       src.ready
		.src_valid          (id_router_011_src_valid),                                                            //          .valid
		.src_data           (id_router_011_src_data),                                                             //          .data
		.src_channel        (id_router_011_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                       //          .endofpacket
	);

	nios_sys_id_router_002 id_router_012 (
		.sink_ready         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ntrreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                            //       src.ready
		.src_valid          (id_router_012_src_valid),                                                            //          .valid
		.src_data           (id_router_012_src_data),                                                             //          .data
		.src_channel        (id_router_012_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                                       //          .endofpacket
	);

	nios_sys_id_router_002 id_router_013 (
		.sink_ready         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (emptyreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                      //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                              //       src.ready
		.src_valid          (id_router_013_src_valid),                                                              //          .valid
		.src_data           (id_router_013_src_data),                                                               //          .data
		.src_channel        (id_router_013_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                                         //          .endofpacket
	);

	nios_sys_id_router_002 id_router_014 (
		.sink_ready         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (emptyreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                      //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                              //       src.ready
		.src_valid          (id_router_014_src_valid),                                                              //          .valid
		.src_data           (id_router_014_src_data),                                                               //          .data
		.src_channel        (id_router_014_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                         //          .endofpacket
	);

	nios_sys_id_router_002 id_router_015 (
		.sink_ready         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (endtsetreg_1_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                        //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                                //       src.ready
		.src_valid          (id_router_015_src_valid),                                                                //          .valid
		.src_data           (id_router_015_src_data),                                                                 //          .data
		.src_channel        (id_router_015_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                           //          .endofpacket
	);

	nios_sys_id_router_002 id_router_016 (
		.sink_ready         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (baseqaddr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                               //       src.ready
		.src_valid          (id_router_016_src_valid),                                                               //          .valid
		.src_data           (id_router_016_src_data),                                                                //          .data
		.src_channel        (id_router_016_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                          //          .endofpacket
	);

	nios_sys_id_router_002 id_router_017 (
		.sink_ready         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (skipaddrreg_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                         //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_017_src_valid),                                                                 //          .valid
		.src_data           (id_router_017_src_data),                                                                  //          .data
		.src_channel        (id_router_017_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                            //          .endofpacket
	);

	nios_sys_id_router_002 id_router_018 (
		.sink_ready         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (knnclasscore_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                        //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                                //       src.ready
		.src_valid          (id_router_018_src_valid),                                                                //          .valid
		.src_data           (id_router_018_src_data),                                                                 //          .data
		.src_channel        (id_router_018_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                           //          .endofpacket
	);

	nios_sys_id_router_002 id_router_019 (
		.sink_ready         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (emptyreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                      //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                              //       src.ready
		.src_valid          (id_router_019_src_valid),                                                              //          .valid
		.src_data           (id_router_019_src_data),                                                               //          .data
		.src_channel        (id_router_019_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                                         //          .endofpacket
	);

	nios_sys_id_router_002 id_router_020 (
		.sink_ready         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (endtsetreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                        //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                                //       src.ready
		.src_valid          (id_router_020_src_valid),                                                                //          .valid
		.src_data           (id_router_020_src_data),                                                                 //          .data
		.src_channel        (id_router_020_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                                           //          .endofpacket
	);

	nios_sys_id_router_002 id_router_021 (
		.sink_ready         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fullreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                     //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                                             //       src.ready
		.src_valid          (id_router_021_src_valid),                                                             //          .valid
		.src_data           (id_router_021_src_data),                                                              //          .data
		.src_channel        (id_router_021_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                                        //          .endofpacket
	);

	nios_sys_id_router_002 id_router_022 (
		.sink_ready         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ntrreg_2_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                    //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_022_src_ready),                                                            //       src.ready
		.src_valid          (id_router_022_src_valid),                                                            //          .valid
		.src_data           (id_router_022_src_data),                                                             //          .data
		.src_channel        (id_router_022_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_022_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_022_src_endofpacket)                                                       //          .endofpacket
	);

	nios_sys_addr_router_003 addr_router_003 (
		.sink_ready         (dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                    //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                    //          .valid
		.src_data           (addr_router_003_src_data),                                                     //          .data
		.src_channel        (addr_router_003_src_channel),                                                  //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                               //          .endofpacket
	);

	nios_sys_addr_router_004 addr_router_004 (
		.sink_ready         (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (distancecore_2_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                                //          .valid
		.src_data           (addr_router_004_src_data),                                                                 //          .data
		.src_channel        (addr_router_004_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                           //          .endofpacket
	);

	nios_sys_addr_router_005 addr_router_005 (
		.sink_ready         (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (distancecore_1_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                                //          .valid
		.src_data           (addr_router_005_src_data),                                                                 //          .data
		.src_channel        (addr_router_005_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                           //          .endofpacket
	);

	nios_sys_addr_router_006 addr_router_006 (
		.sink_ready         (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (distancecore_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                          //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                                //          .valid
		.src_data           (addr_router_006_src_data),                                                                 //          .data
		.src_channel        (addr_router_006_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                                           //          .endofpacket
	);

	nios_sys_id_router_023 id_router_023 (
		.sink_ready         (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cache_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_023_src_ready),                                               //       src.ready
		.src_valid          (id_router_023_src_valid),                                               //          .valid
		.src_data           (id_router_023_src_data),                                                //          .data
		.src_channel        (id_router_023_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_023_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_023_src_endofpacket)                                          //          .endofpacket
	);

	nios_sys_id_router_024 id_router_024 (
		.sink_ready         (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cache_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_024_src_ready),                                               //       src.ready
		.src_valid          (id_router_024_src_valid),                                               //          .valid
		.src_data           (id_router_024_src_data),                                                //          .data
		.src_channel        (id_router_024_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_024_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_024_src_endofpacket)                                          //          .endofpacket
	);

	nios_sys_id_router_025 id_router_025 (
		.sink_ready         (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cache_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_025_src_ready),                                               //       src.ready
		.src_valid          (id_router_025_src_valid),                                               //          .valid
		.src_data           (id_router_025_src_data),                                                //          .data
		.src_channel        (id_router_025_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_025_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_025_src_endofpacket)                                          //          .endofpacket
	);

	nios_sys_addr_router_007 addr_router_007 (
		.sink_ready         (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (distancecore_0_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                                  //          .valid
		.src_data           (addr_router_007_src_data),                                                                   //          .data
		.src_channel        (addr_router_007_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                                             //          .endofpacket
	);

	nios_sys_id_router_026 id_router_026 (
		.sink_ready         (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cache_0_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_026_src_ready),                                               //       src.ready
		.src_valid          (id_router_026_src_valid),                                               //          .valid
		.src_data           (id_router_026_src_data),                                                //          .data
		.src_channel        (id_router_026_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_026_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_026_src_endofpacket)                                          //          .endofpacket
	);

	nios_sys_addr_router_008 addr_router_008 (
		.sink_ready         (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (distancecore_1_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (addr_router_008_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_008_src_valid),                                                                  //          .valid
		.src_data           (addr_router_008_src_data),                                                                   //          .data
		.src_channel        (addr_router_008_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_008_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_008_src_endofpacket)                                                             //          .endofpacket
	);

	nios_sys_id_router_026 id_router_027 (
		.sink_ready         (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cache_1_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_027_src_ready),                                               //       src.ready
		.src_valid          (id_router_027_src_valid),                                               //          .valid
		.src_data           (id_router_027_src_data),                                                //          .data
		.src_channel        (id_router_027_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_027_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_027_src_endofpacket)                                          //          .endofpacket
	);

	nios_sys_addr_router_009 addr_router_009 (
		.sink_ready         (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (distancecore_2_avalon_master_1_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_1_c0_clk),                                                                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (addr_router_009_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_009_src_valid),                                                                  //          .valid
		.src_data           (addr_router_009_src_data),                                                                   //          .data
		.src_channel        (addr_router_009_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_009_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_009_src_endofpacket)                                                             //          .endofpacket
	);

	nios_sys_id_router_026 id_router_028 (
		.sink_ready         (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cache_2_s2_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c2_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_028_src_ready),                                               //       src.ready
		.src_valid          (id_router_028_src_valid),                                               //          .valid
		.src_data           (id_router_028_src_data),                                                //          .data
		.src_channel        (id_router_028_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_028_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_028_src_endofpacket)                                          //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (43),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (63),
		.PKT_BYTE_CNT_H            (52),
		.PKT_BYTE_CNT_L            (50),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (53),
		.PKT_TRANS_COMPRESSED_READ (44),
		.PKT_TRANS_WRITE           (46),
		.PKT_TRANS_READ            (47),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (85),
		.ST_CHANNEL_W              (23),
		.OUT_BYTE_CNT_H            (51),
		.OUT_BURSTWRAP_H           (55),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (7),
		.BURSTWRAP_CONST_VALUE     (7)
	) burst_adapter (
		.clk                   (altpll_0_c0_clk),                     //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                       // reset_in0.reset
		.clk        (altpll_0_c2_clk),                //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.clk        (altpll_0_c0_clk),                    //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.clk        (clk_0),                              //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.clk        (altpll_1_c0_clk),                    //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.clk        (clk_1_clk_in_clk),                   //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_sys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (altpll_0_c2_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (altpll_0_c2_clk),                        //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket),   //          .endofpacket
		.src22_ready         (cmd_xbar_demux_001_src22_ready),         //     src22.ready
		.src22_valid         (cmd_xbar_demux_001_src22_valid),         //          .valid
		.src22_data          (cmd_xbar_demux_001_src22_data),          //          .data
		.src22_channel       (cmd_xbar_demux_001_src22_channel),       //          .channel
		.src22_startofpacket (cmd_xbar_demux_001_src22_startofpacket), //          .startofpacket
		.src22_endofpacket   (cmd_xbar_demux_001_src22_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (altpll_0_c2_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (altpll_0_c2_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (altpll_0_c2_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src5_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux rsp_xbar_demux (
		.clk                (altpll_0_c2_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux rsp_xbar_demux_001 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux rsp_xbar_demux_005 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_011 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_012 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_013 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_014 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_015 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_016 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_017 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_018 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_019 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_020 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_021 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_002 rsp_xbar_demux_022 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_022_src_ready),               //      sink.ready
		.sink_channel       (id_router_022_src_channel),             //          .channel
		.sink_data          (id_router_022_src_data),                //          .data
		.sink_startofpacket (id_router_022_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_022_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_022_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_022_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_022_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_022_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_022_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_022_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_022_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (altpll_0_c2_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (altpll_0_c2_clk),                       //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (crosser_017_out_ready),                 //     sink4.ready
		.sink4_valid          (crosser_017_out_valid),                 //          .valid
		.sink4_channel        (crosser_017_out_channel),               //          .channel
		.sink4_data           (crosser_017_out_data),                  //          .data
		.sink4_startofpacket  (crosser_017_out_startofpacket),         //          .startofpacket
		.sink4_endofpacket    (crosser_017_out_endofpacket),           //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (crosser_018_out_ready),                 //     sink7.ready
		.sink7_valid          (crosser_018_out_valid),                 //          .valid
		.sink7_channel        (crosser_018_out_channel),               //          .channel
		.sink7_data           (crosser_018_out_data),                  //          .data
		.sink7_startofpacket  (crosser_018_out_startofpacket),         //          .startofpacket
		.sink7_endofpacket    (crosser_018_out_endofpacket),           //          .endofpacket
		.sink8_ready          (crosser_019_out_ready),                 //     sink8.ready
		.sink8_valid          (crosser_019_out_valid),                 //          .valid
		.sink8_channel        (crosser_019_out_channel),               //          .channel
		.sink8_data           (crosser_019_out_data),                  //          .data
		.sink8_startofpacket  (crosser_019_out_startofpacket),         //          .startofpacket
		.sink8_endofpacket    (crosser_019_out_endofpacket),           //          .endofpacket
		.sink9_ready          (crosser_020_out_ready),                 //     sink9.ready
		.sink9_valid          (crosser_020_out_valid),                 //          .valid
		.sink9_channel        (crosser_020_out_channel),               //          .channel
		.sink9_data           (crosser_020_out_data),                  //          .data
		.sink9_startofpacket  (crosser_020_out_startofpacket),         //          .startofpacket
		.sink9_endofpacket    (crosser_020_out_endofpacket),           //          .endofpacket
		.sink10_ready         (crosser_021_out_ready),                 //    sink10.ready
		.sink10_valid         (crosser_021_out_valid),                 //          .valid
		.sink10_channel       (crosser_021_out_channel),               //          .channel
		.sink10_data          (crosser_021_out_data),                  //          .data
		.sink10_startofpacket (crosser_021_out_startofpacket),         //          .startofpacket
		.sink10_endofpacket   (crosser_021_out_endofpacket),           //          .endofpacket
		.sink11_ready         (crosser_022_out_ready),                 //    sink11.ready
		.sink11_valid         (crosser_022_out_valid),                 //          .valid
		.sink11_channel       (crosser_022_out_channel),               //          .channel
		.sink11_data          (crosser_022_out_data),                  //          .data
		.sink11_startofpacket (crosser_022_out_startofpacket),         //          .startofpacket
		.sink11_endofpacket   (crosser_022_out_endofpacket),           //          .endofpacket
		.sink12_ready         (crosser_023_out_ready),                 //    sink12.ready
		.sink12_valid         (crosser_023_out_valid),                 //          .valid
		.sink12_channel       (crosser_023_out_channel),               //          .channel
		.sink12_data          (crosser_023_out_data),                  //          .data
		.sink12_startofpacket (crosser_023_out_startofpacket),         //          .startofpacket
		.sink12_endofpacket   (crosser_023_out_endofpacket),           //          .endofpacket
		.sink13_ready         (crosser_024_out_ready),                 //    sink13.ready
		.sink13_valid         (crosser_024_out_valid),                 //          .valid
		.sink13_channel       (crosser_024_out_channel),               //          .channel
		.sink13_data          (crosser_024_out_data),                  //          .data
		.sink13_startofpacket (crosser_024_out_startofpacket),         //          .startofpacket
		.sink13_endofpacket   (crosser_024_out_endofpacket),           //          .endofpacket
		.sink14_ready         (crosser_025_out_ready),                 //    sink14.ready
		.sink14_valid         (crosser_025_out_valid),                 //          .valid
		.sink14_channel       (crosser_025_out_channel),               //          .channel
		.sink14_data          (crosser_025_out_data),                  //          .data
		.sink14_startofpacket (crosser_025_out_startofpacket),         //          .startofpacket
		.sink14_endofpacket   (crosser_025_out_endofpacket),           //          .endofpacket
		.sink15_ready         (crosser_026_out_ready),                 //    sink15.ready
		.sink15_valid         (crosser_026_out_valid),                 //          .valid
		.sink15_channel       (crosser_026_out_channel),               //          .channel
		.sink15_data          (crosser_026_out_data),                  //          .data
		.sink15_startofpacket (crosser_026_out_startofpacket),         //          .startofpacket
		.sink15_endofpacket   (crosser_026_out_endofpacket),           //          .endofpacket
		.sink16_ready         (crosser_027_out_ready),                 //    sink16.ready
		.sink16_valid         (crosser_027_out_valid),                 //          .valid
		.sink16_channel       (crosser_027_out_channel),               //          .channel
		.sink16_data          (crosser_027_out_data),                  //          .data
		.sink16_startofpacket (crosser_027_out_startofpacket),         //          .startofpacket
		.sink16_endofpacket   (crosser_027_out_endofpacket),           //          .endofpacket
		.sink17_ready         (crosser_028_out_ready),                 //    sink17.ready
		.sink17_valid         (crosser_028_out_valid),                 //          .valid
		.sink17_channel       (crosser_028_out_channel),               //          .channel
		.sink17_data          (crosser_028_out_data),                  //          .data
		.sink17_startofpacket (crosser_028_out_startofpacket),         //          .startofpacket
		.sink17_endofpacket   (crosser_028_out_endofpacket),           //          .endofpacket
		.sink18_ready         (crosser_029_out_ready),                 //    sink18.ready
		.sink18_valid         (crosser_029_out_valid),                 //          .valid
		.sink18_channel       (crosser_029_out_channel),               //          .channel
		.sink18_data          (crosser_029_out_data),                  //          .data
		.sink18_startofpacket (crosser_029_out_startofpacket),         //          .startofpacket
		.sink18_endofpacket   (crosser_029_out_endofpacket),           //          .endofpacket
		.sink19_ready         (crosser_030_out_ready),                 //    sink19.ready
		.sink19_valid         (crosser_030_out_valid),                 //          .valid
		.sink19_channel       (crosser_030_out_channel),               //          .channel
		.sink19_data          (crosser_030_out_data),                  //          .data
		.sink19_startofpacket (crosser_030_out_startofpacket),         //          .startofpacket
		.sink19_endofpacket   (crosser_030_out_endofpacket),           //          .endofpacket
		.sink20_ready         (crosser_031_out_ready),                 //    sink20.ready
		.sink20_valid         (crosser_031_out_valid),                 //          .valid
		.sink20_channel       (crosser_031_out_channel),               //          .channel
		.sink20_data          (crosser_031_out_data),                  //          .data
		.sink20_startofpacket (crosser_031_out_startofpacket),         //          .startofpacket
		.sink20_endofpacket   (crosser_031_out_endofpacket),           //          .endofpacket
		.sink21_ready         (crosser_032_out_ready),                 //    sink21.ready
		.sink21_valid         (crosser_032_out_valid),                 //          .valid
		.sink21_channel       (crosser_032_out_channel),               //          .channel
		.sink21_data          (crosser_032_out_data),                  //          .data
		.sink21_startofpacket (crosser_032_out_startofpacket),         //          .startofpacket
		.sink21_endofpacket   (crosser_032_out_endofpacket),           //          .endofpacket
		.sink22_ready         (crosser_033_out_ready),                 //    sink22.ready
		.sink22_valid         (crosser_033_out_valid),                 //          .valid
		.sink22_channel       (crosser_033_out_channel),               //          .channel
		.sink22_data          (crosser_033_out_data),                  //          .data
		.sink22_startofpacket (crosser_033_out_startofpacket),         //          .startofpacket
		.sink22_endofpacket   (crosser_033_out_endofpacket)            //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_003_src2_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_004 cmd_xbar_demux_005 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_004 cmd_xbar_demux_006 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_006_src_ready),             //      sink.ready
		.sink_channel       (addr_router_006_src_channel),           //          .channel
		.sink_data          (addr_router_006_src_data),              //          .data
		.sink_startofpacket (addr_router_006_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_006_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_006_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux_023 cmd_xbar_mux_023 (
		.clk                 (altpll_0_c2_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_023_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_023_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_023_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_023_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_023_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_023_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src0_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_036_out_ready),                 //     sink1.ready
		.sink1_valid         (crosser_036_out_valid),                 //          .valid
		.sink1_channel       (crosser_036_out_channel),               //          .channel
		.sink1_data          (crosser_036_out_data),                  //          .data
		.sink1_startofpacket (crosser_036_out_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (crosser_036_out_endofpacket)            //          .endofpacket
	);

	nios_sys_cmd_xbar_mux_023 cmd_xbar_mux_024 (
		.clk                 (altpll_0_c2_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_024_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_024_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_024_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_024_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_024_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_024_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src1_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src1_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src1_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src1_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_035_out_ready),                 //     sink1.ready
		.sink1_valid         (crosser_035_out_valid),                 //          .valid
		.sink1_channel       (crosser_035_out_channel),               //          .channel
		.sink1_data          (crosser_035_out_data),                  //          .data
		.sink1_startofpacket (crosser_035_out_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (crosser_035_out_endofpacket)            //          .endofpacket
	);

	nios_sys_cmd_xbar_mux_023 cmd_xbar_mux_025 (
		.clk                 (altpll_0_c2_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_025_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_025_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_025_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_025_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_025_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_025_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src2_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src2_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src2_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src2_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (crosser_034_out_ready),                 //     sink1.ready
		.sink1_valid         (crosser_034_out_valid),                 //          .valid
		.sink1_channel       (crosser_034_out_channel),               //          .channel
		.sink1_data          (crosser_034_out_data),                  //          .data
		.sink1_startofpacket (crosser_034_out_startofpacket),         //          .startofpacket
		.sink1_endofpacket   (crosser_034_out_endofpacket)            //          .endofpacket
	);

	nios_sys_rsp_xbar_demux_023 rsp_xbar_demux_023 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_023_src_ready),               //      sink.ready
		.sink_channel       (id_router_023_src_channel),             //          .channel
		.sink_data          (id_router_023_src_data),                //          .data
		.sink_startofpacket (id_router_023_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_023_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_023_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_023_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_023_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_023_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_023_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_023_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_023_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_023_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux_023 rsp_xbar_demux_024 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_024_src_ready),               //      sink.ready
		.sink_channel       (id_router_024_src_channel),             //          .channel
		.sink_data          (id_router_024_src_data),                //          .data
		.sink_startofpacket (id_router_024_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_024_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_024_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_024_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_024_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_024_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_024_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_024_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_024_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_024_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux_023 rsp_xbar_demux_025 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_025_src_ready),               //      sink.ready
		.sink_channel       (id_router_025_src_channel),             //          .channel
		.sink_data          (id_router_025_src_data),                //          .data
		.sink_startofpacket (id_router_025_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_025_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_025_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_025_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_025_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_025_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_025_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_025_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_025_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_025_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_025_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_mux_003 rsp_xbar_mux_003 (
		.clk                 (altpll_0_c2_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_023_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_023_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_023_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_023_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_023_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_023_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_024_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_024_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_024_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_024_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_024_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_024_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_025_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_025_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_025_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_025_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_025_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_025_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_007 cmd_xbar_demux_007 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_007_src_ready),             //      sink.ready
		.sink_channel       (addr_router_007_src_channel),           //          .channel
		.sink_data          (addr_router_007_src_data),              //          .data
		.sink_startofpacket (addr_router_007_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_007_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_007_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_007 rsp_xbar_demux_026 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_026_src_ready),               //      sink.ready
		.sink_channel       (id_router_026_src_channel),             //          .channel
		.sink_data          (id_router_026_src_data),                //          .data
		.sink_startofpacket (id_router_026_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_026_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_026_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_026_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_026_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_026_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_026_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_026_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_026_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_007 cmd_xbar_demux_008 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_008_src_ready),             //      sink.ready
		.sink_channel       (addr_router_008_src_channel),           //          .channel
		.sink_data          (addr_router_008_src_data),              //          .data
		.sink_startofpacket (addr_router_008_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_008_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_008_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_007 rsp_xbar_demux_027 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_027_src_ready),               //      sink.ready
		.sink_channel       (id_router_027_src_channel),             //          .channel
		.sink_data          (id_router_027_src_data),                //          .data
		.sink_startofpacket (id_router_027_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_027_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_027_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_027_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_027_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_027_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_027_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_027_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_027_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_007 cmd_xbar_demux_009 (
		.clk                (altpll_1_c0_clk),                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_009_src_ready),             //      sink.ready
		.sink_channel       (addr_router_009_src_channel),           //          .channel
		.sink_data          (addr_router_009_src_data),              //          .data
		.sink_startofpacket (addr_router_009_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_009_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_009_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux_007 rsp_xbar_demux_028 (
		.clk                (altpll_0_c2_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_028_src_ready),               //      sink.ready
		.sink_channel       (id_router_028_src_channel),             //          .channel
		.sink_data          (id_router_028_src_data),                //          .data
		.sink_startofpacket (id_router_028_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_028_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_028_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_028_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_028_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_028_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_028_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_028_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_028_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (61),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (70),
		.IN_PKT_BYTE_CNT_L             (68),
		.IN_PKT_TRANS_COMPRESSED_READ  (62),
		.IN_PKT_BURSTWRAP_H            (73),
		.IN_PKT_BURSTWRAP_L            (71),
		.IN_PKT_BURST_SIZE_H           (76),
		.IN_PKT_BURST_SIZE_L           (74),
		.IN_PKT_RESPONSE_STATUS_H      (102),
		.IN_PKT_RESPONSE_STATUS_L      (101),
		.IN_PKT_TRANS_EXCLUSIVE        (67),
		.IN_PKT_BURST_TYPE_H           (78),
		.IN_PKT_BURST_TYPE_L           (77),
		.IN_ST_DATA_W                  (103),
		.OUT_PKT_ADDR_H                (43),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (52),
		.OUT_PKT_BYTE_CNT_L            (50),
		.OUT_PKT_TRANS_COMPRESSED_READ (44),
		.OUT_PKT_BURST_SIZE_H          (58),
		.OUT_PKT_BURST_SIZE_L          (56),
		.OUT_PKT_RESPONSE_STATUS_H     (84),
		.OUT_PKT_RESPONSE_STATUS_L     (83),
		.OUT_PKT_TRANS_EXCLUSIVE       (49),
		.OUT_PKT_BURST_TYPE_H          (60),
		.OUT_PKT_BURST_TYPE_L          (59),
		.OUT_ST_DATA_W                 (85),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (altpll_0_c0_clk),                    //       clk.clk
		.reset                (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid             (crosser_out_valid),                  //      sink.valid
		.in_channel           (crosser_out_channel),                //          .channel
		.in_startofpacket     (crosser_out_startofpacket),          //          .startofpacket
		.in_endofpacket       (crosser_out_endofpacket),            //          .endofpacket
		.in_ready             (crosser_out_ready),                  //          .ready
		.in_data              (crosser_out_data),                   //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (43),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (52),
		.IN_PKT_BYTE_CNT_L             (50),
		.IN_PKT_TRANS_COMPRESSED_READ  (44),
		.IN_PKT_BURSTWRAP_H            (55),
		.IN_PKT_BURSTWRAP_L            (53),
		.IN_PKT_BURST_SIZE_H           (58),
		.IN_PKT_BURST_SIZE_L           (56),
		.IN_PKT_RESPONSE_STATUS_H      (84),
		.IN_PKT_RESPONSE_STATUS_L      (83),
		.IN_PKT_TRANS_EXCLUSIVE        (49),
		.IN_PKT_BURST_TYPE_H           (60),
		.IN_PKT_BURST_TYPE_L           (59),
		.IN_ST_DATA_W                  (85),
		.OUT_PKT_ADDR_H                (61),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (70),
		.OUT_PKT_BYTE_CNT_L            (68),
		.OUT_PKT_TRANS_COMPRESSED_READ (62),
		.OUT_PKT_BURST_SIZE_H          (76),
		.OUT_PKT_BURST_SIZE_L          (74),
		.OUT_PKT_RESPONSE_STATUS_H     (102),
		.OUT_PKT_RESPONSE_STATUS_L     (101),
		.OUT_PKT_TRANS_EXCLUSIVE       (67),
		.OUT_PKT_BURST_TYPE_H          (78),
		.OUT_PKT_BURST_TYPE_L          (77),
		.OUT_ST_DATA_W                 (103),
		.ST_CHANNEL_W                  (23),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (altpll_0_c0_clk),                     //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_004_src_valid),             //      sink.valid
		.in_channel           (id_router_004_src_channel),           //          .channel
		.in_startofpacket     (id_router_004_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_004_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_004_src_ready),             //          .ready
		.in_data              (id_router_004_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src4_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src4_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src4_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src4_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src4_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src7_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src7_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src7_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src7_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src7_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src8_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src8_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src8_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src8_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src8_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src9_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src9_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src9_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src9_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src9_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src10_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src10_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src10_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src10_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src10_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src10_data),          //              .data
		.out_ready         (crosser_004_out_ready),                  //           out.ready
		.out_valid         (crosser_004_out_valid),                  //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_004_out_channel),                //              .channel
		.out_data          (crosser_004_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src11_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src11_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src11_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src11_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src11_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src11_data),          //              .data
		.out_ready         (crosser_005_out_ready),                  //           out.ready
		.out_valid         (crosser_005_out_valid),                  //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_005_out_channel),                //              .channel
		.out_data          (crosser_005_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src12_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src12_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src12_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src12_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src12_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src12_data),          //              .data
		.out_ready         (crosser_006_out_ready),                  //           out.ready
		.out_valid         (crosser_006_out_valid),                  //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_006_out_channel),                //              .channel
		.out_data          (crosser_006_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src13_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src13_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src13_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src13_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src13_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src13_data),          //              .data
		.out_ready         (crosser_007_out_ready),                  //           out.ready
		.out_valid         (crosser_007_out_valid),                  //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_007_out_channel),                //              .channel
		.out_data          (crosser_007_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_008 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src14_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src14_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src14_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src14_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src14_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src14_data),          //              .data
		.out_ready         (crosser_008_out_ready),                  //           out.ready
		.out_valid         (crosser_008_out_valid),                  //              .valid
		.out_startofpacket (crosser_008_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_008_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_008_out_channel),                //              .channel
		.out_data          (crosser_008_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_009 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src15_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src15_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src15_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src15_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src15_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src15_data),          //              .data
		.out_ready         (crosser_009_out_ready),                  //           out.ready
		.out_valid         (crosser_009_out_valid),                  //              .valid
		.out_startofpacket (crosser_009_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_009_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_009_out_channel),                //              .channel
		.out_data          (crosser_009_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_010 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src16_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src16_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src16_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src16_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src16_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src16_data),          //              .data
		.out_ready         (crosser_010_out_ready),                  //           out.ready
		.out_valid         (crosser_010_out_valid),                  //              .valid
		.out_startofpacket (crosser_010_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_010_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_010_out_channel),                //              .channel
		.out_data          (crosser_010_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_011 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src17_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src17_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src17_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src17_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src17_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src17_data),          //              .data
		.out_ready         (crosser_011_out_ready),                  //           out.ready
		.out_valid         (crosser_011_out_valid),                  //              .valid
		.out_startofpacket (crosser_011_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_011_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_011_out_channel),                //              .channel
		.out_data          (crosser_011_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_012 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src18_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src18_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src18_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src18_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src18_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src18_data),          //              .data
		.out_ready         (crosser_012_out_ready),                  //           out.ready
		.out_valid         (crosser_012_out_valid),                  //              .valid
		.out_startofpacket (crosser_012_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_012_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_012_out_channel),                //              .channel
		.out_data          (crosser_012_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_013 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src19_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src19_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src19_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src19_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src19_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src19_data),          //              .data
		.out_ready         (crosser_013_out_ready),                  //           out.ready
		.out_valid         (crosser_013_out_valid),                  //              .valid
		.out_startofpacket (crosser_013_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_013_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_013_out_channel),                //              .channel
		.out_data          (crosser_013_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_014 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src20_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src20_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src20_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src20_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src20_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src20_data),          //              .data
		.out_ready         (crosser_014_out_ready),                  //           out.ready
		.out_valid         (crosser_014_out_valid),                  //              .valid
		.out_startofpacket (crosser_014_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_014_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_014_out_channel),                //              .channel
		.out_data          (crosser_014_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_015 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src21_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src21_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src21_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src21_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src21_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src21_data),          //              .data
		.out_ready         (crosser_015_out_ready),                  //           out.ready
		.out_valid         (crosser_015_out_valid),                  //              .valid
		.out_startofpacket (crosser_015_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_015_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_015_out_channel),                //              .channel
		.out_data          (crosser_015_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_016 (
		.in_clk            (altpll_0_c2_clk),                        //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),         //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                        //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),     // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src22_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src22_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src22_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src22_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src22_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src22_data),          //              .data
		.out_ready         (crosser_016_out_ready),                  //           out.ready
		.out_valid         (crosser_016_out_valid),                  //              .valid
		.out_startofpacket (crosser_016_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_016_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_016_out_channel),                //              .channel
		.out_data          (crosser_016_out_data),                   //              .data
		.in_empty          (1'b0),                                   //   (terminated)
		.in_error          (1'b0),                                   //   (terminated)
		.out_empty         (),                                       //   (terminated)
		.out_error         ()                                        //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_017 (
		.in_clk            (altpll_0_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_017_out_ready),                 //           out.ready
		.out_valid         (crosser_017_out_valid),                 //              .valid
		.out_startofpacket (crosser_017_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_017_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_017_out_channel),               //              .channel
		.out_data          (crosser_017_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_018 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_007_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_007_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_007_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_007_src0_data),          //              .data
		.out_ready         (crosser_018_out_ready),                 //           out.ready
		.out_valid         (crosser_018_out_valid),                 //              .valid
		.out_startofpacket (crosser_018_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_018_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_018_out_channel),               //              .channel
		.out_data          (crosser_018_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_019 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_008_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_008_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_008_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_008_src0_data),          //              .data
		.out_ready         (crosser_019_out_ready),                 //           out.ready
		.out_valid         (crosser_019_out_valid),                 //              .valid
		.out_startofpacket (crosser_019_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_019_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_019_out_channel),               //              .channel
		.out_data          (crosser_019_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_020 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_009_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_009_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_009_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_009_src0_data),          //              .data
		.out_ready         (crosser_020_out_ready),                 //           out.ready
		.out_valid         (crosser_020_out_valid),                 //              .valid
		.out_startofpacket (crosser_020_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_020_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_020_out_channel),               //              .channel
		.out_data          (crosser_020_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_021 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_010_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_010_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_010_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_010_src0_data),          //              .data
		.out_ready         (crosser_021_out_ready),                 //           out.ready
		.out_valid         (crosser_021_out_valid),                 //              .valid
		.out_startofpacket (crosser_021_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_021_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_021_out_channel),               //              .channel
		.out_data          (crosser_021_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_022 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_011_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_011_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_011_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_011_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_011_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_011_src0_data),          //              .data
		.out_ready         (crosser_022_out_ready),                 //           out.ready
		.out_valid         (crosser_022_out_valid),                 //              .valid
		.out_startofpacket (crosser_022_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_022_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_022_out_channel),               //              .channel
		.out_data          (crosser_022_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_023 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_012_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_012_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_012_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_012_src0_data),          //              .data
		.out_ready         (crosser_023_out_ready),                 //           out.ready
		.out_valid         (crosser_023_out_valid),                 //              .valid
		.out_startofpacket (crosser_023_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_023_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_023_out_channel),               //              .channel
		.out_data          (crosser_023_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_024 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_013_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_013_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_013_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_013_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_013_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_013_src0_data),          //              .data
		.out_ready         (crosser_024_out_ready),                 //           out.ready
		.out_valid         (crosser_024_out_valid),                 //              .valid
		.out_startofpacket (crosser_024_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_024_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_024_out_channel),               //              .channel
		.out_data          (crosser_024_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_025 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_014_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_014_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_014_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_014_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_014_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_014_src0_data),          //              .data
		.out_ready         (crosser_025_out_ready),                 //           out.ready
		.out_valid         (crosser_025_out_valid),                 //              .valid
		.out_startofpacket (crosser_025_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_025_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_025_out_channel),               //              .channel
		.out_data          (crosser_025_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_026 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_015_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_015_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_015_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_015_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_015_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_015_src0_data),          //              .data
		.out_ready         (crosser_026_out_ready),                 //           out.ready
		.out_valid         (crosser_026_out_valid),                 //              .valid
		.out_startofpacket (crosser_026_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_026_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_026_out_channel),               //              .channel
		.out_data          (crosser_026_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_027 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_016_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_016_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_016_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_016_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_016_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_016_src0_data),          //              .data
		.out_ready         (crosser_027_out_ready),                 //           out.ready
		.out_valid         (crosser_027_out_valid),                 //              .valid
		.out_startofpacket (crosser_027_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_027_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_027_out_channel),               //              .channel
		.out_data          (crosser_027_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_028 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_017_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_017_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_017_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_017_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_017_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_017_src0_data),          //              .data
		.out_ready         (crosser_028_out_ready),                 //           out.ready
		.out_valid         (crosser_028_out_valid),                 //              .valid
		.out_startofpacket (crosser_028_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_028_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_028_out_channel),               //              .channel
		.out_data          (crosser_028_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_029 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_018_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_018_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_018_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_018_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_018_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_018_src0_data),          //              .data
		.out_ready         (crosser_029_out_ready),                 //           out.ready
		.out_valid         (crosser_029_out_valid),                 //              .valid
		.out_startofpacket (crosser_029_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_029_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_029_out_channel),               //              .channel
		.out_data          (crosser_029_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_030 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_019_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_019_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_019_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_019_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_019_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_019_src0_data),          //              .data
		.out_ready         (crosser_030_out_ready),                 //           out.ready
		.out_valid         (crosser_030_out_valid),                 //              .valid
		.out_startofpacket (crosser_030_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_030_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_030_out_channel),               //              .channel
		.out_data          (crosser_030_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_031 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_020_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_020_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_020_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_020_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_020_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_020_src0_data),          //              .data
		.out_ready         (crosser_031_out_ready),                 //           out.ready
		.out_valid         (crosser_031_out_valid),                 //              .valid
		.out_startofpacket (crosser_031_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_031_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_031_out_channel),               //              .channel
		.out_data          (crosser_031_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_032 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_021_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_021_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_021_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_021_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_021_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_021_src0_data),          //              .data
		.out_ready         (crosser_032_out_ready),                 //           out.ready
		.out_valid         (crosser_032_out_valid),                 //              .valid
		.out_startofpacket (crosser_032_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_032_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_032_out_channel),               //              .channel
		.out_data          (crosser_032_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (103),
		.BITS_PER_SYMBOL     (103),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (23),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_033 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_022_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_022_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_022_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_022_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_022_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_022_src0_data),          //              .data
		.out_ready         (crosser_033_out_ready),                 //           out.ready
		.out_valid         (crosser_033_out_valid),                 //              .valid
		.out_startofpacket (crosser_033_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_033_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_033_out_channel),               //              .channel
		.out_data          (crosser_033_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_034 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_034_out_ready),                 //           out.ready
		.out_valid         (crosser_034_out_valid),                 //              .valid
		.out_startofpacket (crosser_034_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_034_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_034_out_channel),               //              .channel
		.out_data          (crosser_034_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_035 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_005_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_005_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_005_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_005_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_005_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_005_src0_data),          //              .data
		.out_ready         (crosser_035_out_ready),                 //           out.ready
		.out_valid         (crosser_035_out_valid),                 //              .valid
		.out_startofpacket (crosser_035_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_035_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_035_out_channel),               //              .channel
		.out_data          (crosser_035_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_036 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_006_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_006_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_006_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_006_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_006_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_006_src0_data),          //              .data
		.out_ready         (crosser_036_out_ready),                 //           out.ready
		.out_valid         (crosser_036_out_valid),                 //              .valid
		.out_startofpacket (crosser_036_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_036_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_036_out_channel),               //              .channel
		.out_data          (crosser_036_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_037 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_023_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_023_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_023_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_023_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_023_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_023_src1_data),          //              .data
		.out_ready         (crosser_037_out_ready),                 //           out.ready
		.out_valid         (crosser_037_out_valid),                 //              .valid
		.out_startofpacket (crosser_037_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_037_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_037_out_channel),               //              .channel
		.out_data          (crosser_037_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_038 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_024_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_024_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_024_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_024_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_024_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_024_src1_data),          //              .data
		.out_ready         (crosser_038_out_ready),                 //           out.ready
		.out_valid         (crosser_038_out_valid),                 //              .valid
		.out_startofpacket (crosser_038_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_038_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_038_out_channel),               //              .channel
		.out_data          (crosser_038_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (87),
		.BITS_PER_SYMBOL     (87),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (4),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_039 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_025_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_025_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_025_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_025_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_025_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_025_src1_data),          //              .data
		.out_ready         (crosser_039_out_ready),                 //           out.ready
		.out_valid         (crosser_039_out_valid),                 //              .valid
		.out_startofpacket (crosser_039_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_039_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_039_out_channel),               //              .channel
		.out_data          (crosser_039_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_040 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_007_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_007_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_007_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_007_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_007_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_007_src0_data),          //              .data
		.out_ready         (crosser_040_out_ready),                 //           out.ready
		.out_valid         (crosser_040_out_valid),                 //              .valid
		.out_startofpacket (crosser_040_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_040_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_040_out_channel),               //              .channel
		.out_data          (crosser_040_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_041 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_026_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_026_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_026_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_026_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_026_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_026_src0_data),          //              .data
		.out_ready         (crosser_041_out_ready),                 //           out.ready
		.out_valid         (crosser_041_out_valid),                 //              .valid
		.out_startofpacket (crosser_041_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_041_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_041_out_channel),               //              .channel
		.out_data          (crosser_041_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_042 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_008_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_008_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_008_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_008_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_008_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_008_src0_data),          //              .data
		.out_ready         (crosser_042_out_ready),                 //           out.ready
		.out_valid         (crosser_042_out_valid),                 //              .valid
		.out_startofpacket (crosser_042_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_042_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_042_out_channel),               //              .channel
		.out_data          (crosser_042_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_043 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_027_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_027_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_027_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_027_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_027_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_027_src0_data),          //              .data
		.out_ready         (crosser_043_out_ready),                 //           out.ready
		.out_valid         (crosser_043_out_valid),                 //              .valid
		.out_startofpacket (crosser_043_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_043_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_043_out_channel),               //              .channel
		.out_data          (crosser_043_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_044 (
		.in_clk            (altpll_1_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c2_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_009_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_009_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_009_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_009_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_009_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_009_src0_data),          //              .data
		.out_ready         (crosser_044_out_ready),                 //           out.ready
		.out_valid         (crosser_044_out_valid),                 //              .valid
		.out_startofpacket (crosser_044_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_044_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_044_out_channel),               //              .channel
		.out_data          (crosser_044_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (85),
		.BITS_PER_SYMBOL     (85),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_045 (
		.in_clk            (altpll_0_c2_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (altpll_1_c0_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_028_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_028_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_028_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_028_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_028_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_028_src0_data),          //              .data
		.out_ready         (crosser_045_out_ready),                 //           out.ready
		.out_valid         (crosser_045_out_valid),                 //              .valid
		.out_startofpacket (crosser_045_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_045_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_045_out_channel),               //              .channel
		.out_data          (crosser_045_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	nios_sys_irq_mapper irq_mapper (
		.clk           (altpll_0_c2_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

endmodule
