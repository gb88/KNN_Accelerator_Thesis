library ieee; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 
use work.common_types.all;
use ieee.math_real.all;

entity AvInterface is 
	port
	(	
		clk,
		reset_n,
		read,
		write,
		chipselect	: in std_logic;
		address		: in std_logic_vector(4 downto 0);
		readdata	: out std_logic_vector(31 downto 0);
		writedata	: in std_logic_vector(31 downto 0);
		ClOut 		: in std_logic_vector(CLASS_WIDTH-1 downto 0);
		NVot:		in std_logic_vector(INTEGER(ceil(log2(real(MAX_KSET_SIZE)))) downto 0);
		StartCl		: out std_logic;
		KVal:		 out std_logic_vector(K_WIDTH-1 downto 0);
		EndClass	: in std_logic;
		DistIn:			in DistArray(MAX_KSET_SIZE-1 downto 0);
		Overflow:	 in std_logic
	);		
end AvInterface; 

architecture Structural of AvInterface is 	 

begin 
	process(clk, reset_n) 
	begin
		if reset_n = '0' then
			readdata <= (others=>'0');
		elsif(rising_edge(clk)) then
			if(chipselect='1')then
				if(read='1')then
					case address is 
						when "00000" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(0);
						when "00001" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(1);
						when "00010" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(2);
						when "00011" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(3);
						when "00100" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(4);
						when "00101" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(5);
						when "00110" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(6);
						when "00111" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(7);
						when "01000" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(8);
						when "01001" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(9);
						when "01010" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(10);
						when "01011" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(11);
						when "01100" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(12);
						when "01101" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(13);
						when "01110" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(14);
						when "01111" =>
							readdata(31 downto 16) <= (Others => '0');
							readdata(15 downto 0) <= DistIn(15);
						when "10000" =>
							readdata(31 downto CLASS_WIDTH) <= (Others => '0');
							readdata(CLASS_WIDTH-1 downto 0) <= ClOut;
						when "10001" =>
							readdata(31 downto INTEGER(ceil(log2(real(MAX_KSET_SIZE))))+1) <= (Others => '0');
							readdata(INTEGER(ceil(log2(real(MAX_KSET_SIZE)))) downto 0) <= NVot;
						when "10010" =>
							readdata(31 downto 1) <= (Others => '0');
							readdata(0) <= EndClass;
						when "10011" =>
							readdata(31 downto 1) <= (Others =>'0');
							readdata(0) <= Overflow;
						when others =>
							readdata <= (others=>'0');
					end case;
				end if;
				if (write='1') then
					case address is
						when "10100" =>
							KVal <= writedata(K_WIDTH-1 downto 0);
						when "10101" =>
							StartCl <= writedata(0);
						when others =>
					end case;
				end if;
			end if;
		end if;
	end process;
	
end structural;