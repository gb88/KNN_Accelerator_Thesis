library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.EucDisPkg.all;
use work.common_types.all;

entity EucDis is
	port 
	(
		Clk : in std_logic;
		Reset : in std_logic; --si pu� togliere
		DimT : in std_logic_vector(DIM_WIDTH-1 downto 0);
		DimQ : in std_logic_vector(DIM_WIDTH-1 downto 0);
		SumEn: in std_logic;
		SubEn: in std_logic;
		SumReset: in std_logic;
		Overflow: out std_logic;
		Dist: out std_logic_vector(DISTANCE_WIDTH-1 downto 0)
	);
end EucDis;

architecture Structural of EucDis is

	signal OverflowSubDimxS: std_logic;
	signal OverflowSumxS: std_logic;
	signal SubDimxD: std_logic_vector(DIM_WIDTH-1 downto 0);
	signal TwoPowerxD: std_logic_vector(DIM_WIDTH*2-3 downto 0);
	
	begin 
		SubDimBlk : SubDim port map (Clk, DimT, DimQ, SubEn, OverflowSubDimxS, SubDimxD);
		TwoPowerBlk : TwoPower port map (Clk, SubDimxD, TwoPowerxD);
		SummationBlk : Summation port map (Clk, SumReset, SumEn, TwoPowerxD, OverflowSumxS, Dist);
		Overflow <= OverflowSubDimxS or OverflowSumxS;
		
end Structural;